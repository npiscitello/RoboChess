// nios_system.v

// Generated using ACDS version 13.0 156 at 2013.06.06.14:41:08

`timescale 1 ps / 1 ps
module nios_system (
		input  wire        reset_n,                              //                   clk_clk_in_reset.reset_n
		inout  wire [31:0] GPIO_0_to_and_from_the_Expansion_JP1, //   Expansion_JP1_external_interface.export
		output wire [9:0]  LEDG_from_the_Green_LEDs,             //      Green_LEDs_external_interface.export
		output wire [11:0] zs_addr_from_the_sdram,               //                         sdram_wire.addr
		output wire [1:0]  zs_ba_from_the_sdram,                 //                                   .ba
		output wire        zs_cas_n_from_the_sdram,              //                                   .cas_n
		output wire        zs_cke_from_the_sdram,                //                                   .cke
		output wire        zs_cs_n_from_the_sdram,               //                                   .cs_n
		inout  wire [15:0] zs_dq_to_and_from_the_sdram,          //                                   .dq
		output wire [1:0]  zs_dqm_from_the_sdram,                //                                   .dqm
		output wire        zs_ras_n_from_the_sdram,              //                                   .ras_n
		output wire        zs_we_n_from_the_sdram,               //                                   .we_n
		inout  wire [31:0] GPIO_1_to_and_from_the_Expansion_JP2, //   Expansion_JP2_external_interface.export
		input  wire        UART_RXD_to_the_Serial_port,          //     Serial_port_external_interface.RXD
		output wire        UART_TXD_from_the_Serial_port,        //                                   .TXD
		input  wire        clk,                                  //                         clk_clk_in.clk
		input  wire [2:0]  KEY_to_the_Pushbuttons,               //     Pushbuttons_external_interface.export
		input  wire [9:0]  SW_to_the_Slider_switches,            // Slider_switches_external_interface.export
		output wire [7:0]  HEX0_from_the_HEX3_HEX0,              //       HEX3_HEX0_external_interface.HEX0
		output wire [7:0]  HEX1_from_the_HEX3_HEX0,              //                                   .HEX1
		output wire [7:0]  HEX2_from_the_HEX3_HEX0,              //                                   .HEX2
		output wire [7:0]  HEX3_from_the_HEX3_HEX0               //                                   .HEX3
	);

	wire          cpu_instruction_master_waitrequest;                                                                              // cpu_instruction_master_translator:av_waitrequest -> cpu:i_waitrequest
	wire   [27:0] cpu_instruction_master_address;                                                                                  // cpu:i_address -> cpu_instruction_master_translator:av_address
	wire          cpu_instruction_master_read;                                                                                     // cpu:i_read -> cpu_instruction_master_translator:av_read
	wire   [31:0] cpu_instruction_master_readdata;                                                                                 // cpu_instruction_master_translator:av_readdata -> cpu:i_readdata
	wire          cpu_data_master_waitrequest;                                                                                     // cpu_data_master_translator:av_waitrequest -> cpu:d_waitrequest
	wire   [31:0] cpu_data_master_writedata;                                                                                       // cpu:d_writedata -> cpu_data_master_translator:av_writedata
	wire   [28:0] cpu_data_master_address;                                                                                         // cpu:d_address -> cpu_data_master_translator:av_address
	wire          cpu_data_master_write;                                                                                           // cpu:d_write -> cpu_data_master_translator:av_write
	wire          cpu_data_master_read;                                                                                            // cpu:d_read -> cpu_data_master_translator:av_read
	wire   [31:0] cpu_data_master_readdata;                                                                                        // cpu_data_master_translator:av_readdata -> cpu:d_readdata
	wire          cpu_data_master_debugaccess;                                                                                     // cpu:jtag_debug_module_debugaccess_to_roms -> cpu_data_master_translator:av_debugaccess
	wire    [3:0] cpu_data_master_byteenable;                                                                                      // cpu:d_byteenable -> cpu_data_master_translator:av_byteenable
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                                                // cpu:jtag_debug_module_waitrequest -> cpu_jtag_debug_module_translator:av_waitrequest
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                                  // cpu_jtag_debug_module_translator:av_writedata -> cpu:jtag_debug_module_writedata
	wire    [8:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_address;                                                    // cpu_jtag_debug_module_translator:av_address -> cpu:jtag_debug_module_address
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_write;                                                      // cpu_jtag_debug_module_translator:av_write -> cpu:jtag_debug_module_write
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_read;                                                       // cpu_jtag_debug_module_translator:av_read -> cpu:jtag_debug_module_read
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                                   // cpu:jtag_debug_module_readdata -> cpu_jtag_debug_module_translator:av_readdata
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                                // cpu_jtag_debug_module_translator:av_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                                 // cpu_jtag_debug_module_translator:av_byteenable -> cpu:jtag_debug_module_byteenable
	wire   [31:0] onchip_memory_s1_translator_avalon_anti_slave_0_writedata;                                                       // Onchip_memory_s1_translator:av_writedata -> Onchip_memory:writedata
	wire   [10:0] onchip_memory_s1_translator_avalon_anti_slave_0_address;                                                         // Onchip_memory_s1_translator:av_address -> Onchip_memory:address
	wire          onchip_memory_s1_translator_avalon_anti_slave_0_chipselect;                                                      // Onchip_memory_s1_translator:av_chipselect -> Onchip_memory:chipselect
	wire          onchip_memory_s1_translator_avalon_anti_slave_0_clken;                                                           // Onchip_memory_s1_translator:av_clken -> Onchip_memory:clken
	wire          onchip_memory_s1_translator_avalon_anti_slave_0_write;                                                           // Onchip_memory_s1_translator:av_write -> Onchip_memory:write
	wire   [31:0] onchip_memory_s1_translator_avalon_anti_slave_0_readdata;                                                        // Onchip_memory:readdata -> Onchip_memory_s1_translator:av_readdata
	wire    [3:0] onchip_memory_s1_translator_avalon_anti_slave_0_byteenable;                                                      // Onchip_memory_s1_translator:av_byteenable -> Onchip_memory:byteenable
	wire          sdram_s1_translator_avalon_anti_slave_0_waitrequest;                                                             // sdram:za_waitrequest -> sdram_s1_translator:av_waitrequest
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_writedata;                                                               // sdram_s1_translator:av_writedata -> sdram:az_data
	wire   [21:0] sdram_s1_translator_avalon_anti_slave_0_address;                                                                 // sdram_s1_translator:av_address -> sdram:az_addr
	wire          sdram_s1_translator_avalon_anti_slave_0_chipselect;                                                              // sdram_s1_translator:av_chipselect -> sdram:az_cs
	wire          sdram_s1_translator_avalon_anti_slave_0_write;                                                                   // sdram_s1_translator:av_write -> sdram:az_wr_n
	wire          sdram_s1_translator_avalon_anti_slave_0_read;                                                                    // sdram_s1_translator:av_read -> sdram:az_rd_n
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_readdata;                                                                // sdram:za_data -> sdram_s1_translator:av_readdata
	wire          sdram_s1_translator_avalon_anti_slave_0_readdatavalid;                                                           // sdram:za_valid -> sdram_s1_translator:av_readdatavalid
	wire    [1:0] sdram_s1_translator_avalon_anti_slave_0_byteenable;                                                              // sdram_s1_translator:av_byteenable -> sdram:az_be_n
	wire   [31:0] onchip_memory_sram_s1_translator_avalon_anti_slave_0_writedata;                                                  // Onchip_memory_SRAM_s1_translator:av_writedata -> Onchip_memory_SRAM:writedata
	wire   [10:0] onchip_memory_sram_s1_translator_avalon_anti_slave_0_address;                                                    // Onchip_memory_SRAM_s1_translator:av_address -> Onchip_memory_SRAM:address
	wire          onchip_memory_sram_s1_translator_avalon_anti_slave_0_chipselect;                                                 // Onchip_memory_SRAM_s1_translator:av_chipselect -> Onchip_memory_SRAM:chipselect
	wire          onchip_memory_sram_s1_translator_avalon_anti_slave_0_clken;                                                      // Onchip_memory_SRAM_s1_translator:av_clken -> Onchip_memory_SRAM:clken
	wire          onchip_memory_sram_s1_translator_avalon_anti_slave_0_write;                                                      // Onchip_memory_SRAM_s1_translator:av_write -> Onchip_memory_SRAM:write
	wire   [31:0] onchip_memory_sram_s1_translator_avalon_anti_slave_0_readdata;                                                   // Onchip_memory_SRAM:readdata -> Onchip_memory_SRAM_s1_translator:av_readdata
	wire    [3:0] onchip_memory_sram_s1_translator_avalon_anti_slave_0_byteenable;                                                 // Onchip_memory_SRAM_s1_translator:av_byteenable -> Onchip_memory_SRAM:byteenable
	wire   [31:0] onchip_memory_s2_translator_avalon_anti_slave_0_writedata;                                                       // Onchip_memory_s2_translator:av_writedata -> Onchip_memory:writedata2
	wire   [10:0] onchip_memory_s2_translator_avalon_anti_slave_0_address;                                                         // Onchip_memory_s2_translator:av_address -> Onchip_memory:address2
	wire          onchip_memory_s2_translator_avalon_anti_slave_0_chipselect;                                                      // Onchip_memory_s2_translator:av_chipselect -> Onchip_memory:chipselect2
	wire          onchip_memory_s2_translator_avalon_anti_slave_0_clken;                                                           // Onchip_memory_s2_translator:av_clken -> Onchip_memory:clken2
	wire          onchip_memory_s2_translator_avalon_anti_slave_0_write;                                                           // Onchip_memory_s2_translator:av_write -> Onchip_memory:write2
	wire   [31:0] onchip_memory_s2_translator_avalon_anti_slave_0_readdata;                                                        // Onchip_memory:readdata2 -> Onchip_memory_s2_translator:av_readdata
	wire    [3:0] onchip_memory_s2_translator_avalon_anti_slave_0_byteenable;                                                      // Onchip_memory_s2_translator:av_byteenable -> Onchip_memory:byteenable2
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                          // JTAG_UART:av_waitrequest -> JTAG_UART_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                            // JTAG_UART_avalon_jtag_slave_translator:av_writedata -> JTAG_UART:av_writedata
	wire    [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                              // JTAG_UART_avalon_jtag_slave_translator:av_address -> JTAG_UART:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                           // JTAG_UART_avalon_jtag_slave_translator:av_chipselect -> JTAG_UART:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                                // JTAG_UART_avalon_jtag_slave_translator:av_write -> JTAG_UART:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                                 // JTAG_UART_avalon_jtag_slave_translator:av_read -> JTAG_UART:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                             // JTAG_UART:av_readdata -> JTAG_UART_avalon_jtag_slave_translator:av_readdata
	wire   [15:0] interval_timer_s1_translator_avalon_anti_slave_0_writedata;                                                      // Interval_timer_s1_translator:av_writedata -> Interval_timer:writedata
	wire    [2:0] interval_timer_s1_translator_avalon_anti_slave_0_address;                                                        // Interval_timer_s1_translator:av_address -> Interval_timer:address
	wire          interval_timer_s1_translator_avalon_anti_slave_0_chipselect;                                                     // Interval_timer_s1_translator:av_chipselect -> Interval_timer:chipselect
	wire          interval_timer_s1_translator_avalon_anti_slave_0_write;                                                          // Interval_timer_s1_translator:av_write -> Interval_timer:write_n
	wire   [15:0] interval_timer_s1_translator_avalon_anti_slave_0_readdata;                                                       // Interval_timer:readdata -> Interval_timer_s1_translator:av_readdata
	wire    [0:0] sysid_control_slave_translator_avalon_anti_slave_0_address;                                                      // sysid_control_slave_translator:av_address -> sysid:address
	wire   [31:0] sysid_control_slave_translator_avalon_anti_slave_0_readdata;                                                     // sysid:readdata -> sysid_control_slave_translator:av_readdata
	wire   [31:0] green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                                  // Green_LEDs_avalon_parallel_port_slave_translator:av_writedata -> Green_LEDs:writedata
	wire    [1:0] green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                                    // Green_LEDs_avalon_parallel_port_slave_translator:av_address -> Green_LEDs:address
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                                 // Green_LEDs_avalon_parallel_port_slave_translator:av_chipselect -> Green_LEDs:chipselect
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                      // Green_LEDs_avalon_parallel_port_slave_translator:av_write -> Green_LEDs:write
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                       // Green_LEDs_avalon_parallel_port_slave_translator:av_read -> Green_LEDs:read
	wire   [31:0] green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                                   // Green_LEDs:readdata -> Green_LEDs_avalon_parallel_port_slave_translator:av_readdata
	wire    [3:0] green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                                 // Green_LEDs_avalon_parallel_port_slave_translator:av_byteenable -> Green_LEDs:byteenable
	wire   [31:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                                   // HEX3_HEX0_avalon_parallel_port_slave_translator:av_writedata -> HEX3_HEX0:writedata
	wire    [1:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                                     // HEX3_HEX0_avalon_parallel_port_slave_translator:av_address -> HEX3_HEX0:address
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                                  // HEX3_HEX0_avalon_parallel_port_slave_translator:av_chipselect -> HEX3_HEX0:chipselect
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                       // HEX3_HEX0_avalon_parallel_port_slave_translator:av_write -> HEX3_HEX0:write
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                        // HEX3_HEX0_avalon_parallel_port_slave_translator:av_read -> HEX3_HEX0:read
	wire   [31:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                                    // HEX3_HEX0:readdata -> HEX3_HEX0_avalon_parallel_port_slave_translator:av_readdata
	wire    [3:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                                  // HEX3_HEX0_avalon_parallel_port_slave_translator:av_byteenable -> HEX3_HEX0:byteenable
	wire   [31:0] slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                             // Slider_switches_avalon_parallel_port_slave_translator:av_writedata -> Slider_switches:writedata
	wire    [1:0] slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                               // Slider_switches_avalon_parallel_port_slave_translator:av_address -> Slider_switches:address
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                            // Slider_switches_avalon_parallel_port_slave_translator:av_chipselect -> Slider_switches:chipselect
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                 // Slider_switches_avalon_parallel_port_slave_translator:av_write -> Slider_switches:write
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                  // Slider_switches_avalon_parallel_port_slave_translator:av_read -> Slider_switches:read
	wire   [31:0] slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                              // Slider_switches:readdata -> Slider_switches_avalon_parallel_port_slave_translator:av_readdata
	wire    [3:0] slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                            // Slider_switches_avalon_parallel_port_slave_translator:av_byteenable -> Slider_switches:byteenable
	wire   [31:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                                 // Pushbuttons_avalon_parallel_port_slave_translator:av_writedata -> Pushbuttons:writedata
	wire    [1:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                                   // Pushbuttons_avalon_parallel_port_slave_translator:av_address -> Pushbuttons:address
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                                // Pushbuttons_avalon_parallel_port_slave_translator:av_chipselect -> Pushbuttons:chipselect
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                     // Pushbuttons_avalon_parallel_port_slave_translator:av_write -> Pushbuttons:write
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                      // Pushbuttons_avalon_parallel_port_slave_translator:av_read -> Pushbuttons:read
	wire   [31:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                                  // Pushbuttons:readdata -> Pushbuttons_avalon_parallel_port_slave_translator:av_readdata
	wire    [3:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                                // Pushbuttons_avalon_parallel_port_slave_translator:av_byteenable -> Pushbuttons:byteenable
	wire   [31:0] expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                               // Expansion_JP1_avalon_parallel_port_slave_translator:av_writedata -> Expansion_JP1:writedata
	wire    [1:0] expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                                 // Expansion_JP1_avalon_parallel_port_slave_translator:av_address -> Expansion_JP1:address
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                              // Expansion_JP1_avalon_parallel_port_slave_translator:av_chipselect -> Expansion_JP1:chipselect
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                   // Expansion_JP1_avalon_parallel_port_slave_translator:av_write -> Expansion_JP1:write
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                    // Expansion_JP1_avalon_parallel_port_slave_translator:av_read -> Expansion_JP1:read
	wire   [31:0] expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                                // Expansion_JP1:readdata -> Expansion_JP1_avalon_parallel_port_slave_translator:av_readdata
	wire    [3:0] expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                              // Expansion_JP1_avalon_parallel_port_slave_translator:av_byteenable -> Expansion_JP1:byteenable
	wire   [31:0] expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                               // Expansion_JP2_avalon_parallel_port_slave_translator:av_writedata -> Expansion_JP2:writedata
	wire    [1:0] expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                                 // Expansion_JP2_avalon_parallel_port_slave_translator:av_address -> Expansion_JP2:address
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                              // Expansion_JP2_avalon_parallel_port_slave_translator:av_chipselect -> Expansion_JP2:chipselect
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                   // Expansion_JP2_avalon_parallel_port_slave_translator:av_write -> Expansion_JP2:write
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                    // Expansion_JP2_avalon_parallel_port_slave_translator:av_read -> Expansion_JP2:read
	wire   [31:0] expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                                // Expansion_JP2:readdata -> Expansion_JP2_avalon_parallel_port_slave_translator:av_readdata
	wire    [3:0] expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                              // Expansion_JP2_avalon_parallel_port_slave_translator:av_byteenable -> Expansion_JP2:byteenable
	wire   [31:0] serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_writedata;                                         // Serial_port_avalon_rs232_slave_translator:av_writedata -> Serial_port:writedata
	wire    [0:0] serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_address;                                           // Serial_port_avalon_rs232_slave_translator:av_address -> Serial_port:address
	wire          serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_chipselect;                                        // Serial_port_avalon_rs232_slave_translator:av_chipselect -> Serial_port:chipselect
	wire          serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_write;                                             // Serial_port_avalon_rs232_slave_translator:av_write -> Serial_port:write
	wire          serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_read;                                              // Serial_port_avalon_rs232_slave_translator:av_read -> Serial_port:read
	wire   [31:0] serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_readdata;                                          // Serial_port:readdata -> Serial_port_avalon_rs232_slave_translator:av_readdata
	wire    [3:0] serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_byteenable;                                        // Serial_port_avalon_rs232_slave_translator:av_byteenable -> Serial_port:byteenable
	wire   [31:0] onchip_memory_sram_s2_translator_avalon_anti_slave_0_writedata;                                                  // Onchip_memory_SRAM_s2_translator:av_writedata -> Onchip_memory_SRAM:writedata2
	wire   [10:0] onchip_memory_sram_s2_translator_avalon_anti_slave_0_address;                                                    // Onchip_memory_SRAM_s2_translator:av_address -> Onchip_memory_SRAM:address2
	wire          onchip_memory_sram_s2_translator_avalon_anti_slave_0_chipselect;                                                 // Onchip_memory_SRAM_s2_translator:av_chipselect -> Onchip_memory_SRAM:chipselect2
	wire          onchip_memory_sram_s2_translator_avalon_anti_slave_0_clken;                                                      // Onchip_memory_SRAM_s2_translator:av_clken -> Onchip_memory_SRAM:clken2
	wire          onchip_memory_sram_s2_translator_avalon_anti_slave_0_write;                                                      // Onchip_memory_SRAM_s2_translator:av_write -> Onchip_memory_SRAM:write2
	wire   [31:0] onchip_memory_sram_s2_translator_avalon_anti_slave_0_readdata;                                                   // Onchip_memory_SRAM:readdata2 -> Onchip_memory_SRAM_s2_translator:av_readdata
	wire    [3:0] onchip_memory_sram_s2_translator_avalon_anti_slave_0_byteenable;                                                 // Onchip_memory_SRAM_s2_translator:av_byteenable -> Onchip_memory_SRAM:byteenable2
	wire          cpu_instruction_master_translator_avalon_universal_master_0_waitrequest;                                         // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_instruction_master_translator_avalon_universal_master_0_burstcount;                                          // cpu_instruction_master_translator:uav_burstcount -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_writedata;                                           // cpu_instruction_master_translator:uav_writedata -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [28:0] cpu_instruction_master_translator_avalon_universal_master_0_address;                                             // cpu_instruction_master_translator:uav_address -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_instruction_master_translator_avalon_universal_master_0_lock;                                                // cpu_instruction_master_translator:uav_lock -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_instruction_master_translator_avalon_universal_master_0_write;                                               // cpu_instruction_master_translator:uav_write -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_instruction_master_translator_avalon_universal_master_0_read;                                                // cpu_instruction_master_translator:uav_read -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_readdata;                                            // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_instruction_master_translator:uav_readdata
	wire          cpu_instruction_master_translator_avalon_universal_master_0_debugaccess;                                         // cpu_instruction_master_translator:uav_debugaccess -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_instruction_master_translator_avalon_universal_master_0_byteenable;                                          // cpu_instruction_master_translator:uav_byteenable -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid;                                       // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_instruction_master_translator:uav_readdatavalid
	wire          cpu_data_master_translator_avalon_universal_master_0_waitrequest;                                                // cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_data_master_translator_avalon_universal_master_0_burstcount;                                                 // cpu_data_master_translator:uav_burstcount -> cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_writedata;                                                  // cpu_data_master_translator:uav_writedata -> cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [28:0] cpu_data_master_translator_avalon_universal_master_0_address;                                                    // cpu_data_master_translator:uav_address -> cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_data_master_translator_avalon_universal_master_0_lock;                                                       // cpu_data_master_translator:uav_lock -> cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_data_master_translator_avalon_universal_master_0_write;                                                      // cpu_data_master_translator:uav_write -> cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_data_master_translator_avalon_universal_master_0_read;                                                       // cpu_data_master_translator:uav_read -> cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_readdata;                                                   // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_data_master_translator:uav_readdata
	wire          cpu_data_master_translator_avalon_universal_master_0_debugaccess;                                                // cpu_data_master_translator:uav_debugaccess -> cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_data_master_translator_avalon_universal_master_0_byteenable;                                                 // cpu_data_master_translator:uav_byteenable -> cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                                              // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_data_master_translator:uav_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // cpu_jtag_debug_module_translator:uav_waitrequest -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_jtag_debug_module_translator:uav_writedata
	wire   [28:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                                      // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_jtag_debug_module_translator:uav_address
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                                        // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_jtag_debug_module_translator:uav_write
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_jtag_debug_module_translator:uav_lock
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_jtag_debug_module_translator:uav_read
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // cpu_jtag_debug_module_translator:uav_readdata -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // cpu_jtag_debug_module_translator:uav_readdatavalid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_jtag_debug_module_translator:uav_byteenable
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                       // Onchip_memory_s1_translator:uav_waitrequest -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                        // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> Onchip_memory_s1_translator:uav_burstcount
	wire   [31:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                         // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> Onchip_memory_s1_translator:uav_writedata
	wire   [28:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address;                                           // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> Onchip_memory_s1_translator:uav_address
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write;                                             // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> Onchip_memory_s1_translator:uav_write
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                              // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> Onchip_memory_s1_translator:uav_lock
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read;                                              // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> Onchip_memory_s1_translator:uav_read
	wire   [31:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                          // Onchip_memory_s1_translator:uav_readdata -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                     // Onchip_memory_s1_translator:uav_readdatavalid -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                       // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Onchip_memory_s1_translator:uav_debugaccess
	wire    [3:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                        // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> Onchip_memory_s1_translator:uav_byteenable
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                      // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                              // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                       // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                      // Onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                             // Onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                   // Onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                           // Onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                    // Onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                   // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                 // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                  // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                 // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                               // sdram_s1_translator:uav_waitrequest -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                // sdram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_s1_translator:uav_burstcount
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                 // sdram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_s1_translator:uav_writedata
	wire   [28:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                   // sdram_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_s1_translator:uav_address
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                     // sdram_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_s1_translator:uav_write
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                      // sdram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_s1_translator:uav_lock
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                      // sdram_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_s1_translator:uav_read
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                  // sdram_s1_translator:uav_readdata -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                             // sdram_s1_translator:uav_readdatavalid -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                               // sdram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_s1_translator:uav_debugaccess
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                // sdram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_s1_translator:uav_byteenable
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                        // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                              // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                      // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [86:0] sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                               // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                              // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                     // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                           // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                   // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [86:0] sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                            // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                           // sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                         // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [17:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                          // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                         // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                         // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                          // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                         // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // Onchip_memory_SRAM_s1_translator:uav_waitrequest -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> Onchip_memory_SRAM_s1_translator:uav_burstcount
	wire   [31:0] onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> Onchip_memory_SRAM_s1_translator:uav_writedata
	wire   [28:0] onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:m0_address -> Onchip_memory_SRAM_s1_translator:uav_address
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:m0_write -> Onchip_memory_SRAM_s1_translator:uav_write
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:m0_lock -> Onchip_memory_SRAM_s1_translator:uav_lock
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:m0_read -> Onchip_memory_SRAM_s1_translator:uav_read
	wire   [31:0] onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // Onchip_memory_SRAM_s1_translator:uav_readdata -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // Onchip_memory_SRAM_s1_translator:uav_readdatavalid -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Onchip_memory_SRAM_s1_translator:uav_debugaccess
	wire    [3:0] onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> Onchip_memory_SRAM_s1_translator:uav_byteenable
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                       // Onchip_memory_s2_translator:uav_waitrequest -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_burstcount;                                        // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:m0_burstcount -> Onchip_memory_s2_translator:uav_burstcount
	wire   [31:0] onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_writedata;                                         // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:m0_writedata -> Onchip_memory_s2_translator:uav_writedata
	wire   [28:0] onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_address;                                           // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:m0_address -> Onchip_memory_s2_translator:uav_address
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_write;                                             // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:m0_write -> Onchip_memory_s2_translator:uav_write
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_lock;                                              // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:m0_lock -> Onchip_memory_s2_translator:uav_lock
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_read;                                              // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:m0_read -> Onchip_memory_s2_translator:uav_read
	wire   [31:0] onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_readdata;                                          // Onchip_memory_s2_translator:uav_readdata -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                     // Onchip_memory_s2_translator:uav_readdatavalid -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                       // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Onchip_memory_s2_translator:uav_debugaccess
	wire    [3:0] onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_byteenable;                                        // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:m0_byteenable -> Onchip_memory_s2_translator:uav_byteenable
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_valid;                                      // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rf_source_valid -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                              // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] onchip_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_data;                                       // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rf_source_data -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_ready;                                      // Onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                             // Onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                   // Onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                           // Onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                    // Onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                   // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                 // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] onchip_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                  // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                 // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // JTAG_UART_avalon_jtag_slave_translator:uav_waitrequest -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> JTAG_UART_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                              // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> JTAG_UART_avalon_jtag_slave_translator:uav_writedata
	wire   [28:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                                // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> JTAG_UART_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                                  // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> JTAG_UART_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                   // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> JTAG_UART_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                                   // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> JTAG_UART_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                               // JTAG_UART_avalon_jtag_slave_translator:uav_readdata -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // JTAG_UART_avalon_jtag_slave_translator:uav_readdatavalid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> JTAG_UART_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> JTAG_UART_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                            // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // Interval_timer_s1_translator:uav_waitrequest -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> Interval_timer_s1_translator:uav_burstcount
	wire   [31:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> Interval_timer_s1_translator:uav_writedata
	wire   [28:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                          // Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> Interval_timer_s1_translator:uav_address
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                            // Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> Interval_timer_s1_translator:uav_write
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                             // Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> Interval_timer_s1_translator:uav_lock
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                             // Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> Interval_timer_s1_translator:uav_read
	wire   [31:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // Interval_timer_s1_translator:uav_readdata -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // Interval_timer_s1_translator:uav_readdatavalid -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Interval_timer_s1_translator:uav_debugaccess
	wire    [3:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> Interval_timer_s1_translator:uav_byteenable
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // Interval_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // Interval_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // Interval_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	wire   [28:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                                        // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	wire    [3:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                  // Green_LEDs_avalon_parallel_port_slave_translator:uav_waitrequest -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                   // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Green_LEDs_avalon_parallel_port_slave_translator:uav_burstcount
	wire   [31:0] green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                    // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Green_LEDs_avalon_parallel_port_slave_translator:uav_writedata
	wire   [28:0] green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                      // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> Green_LEDs_avalon_parallel_port_slave_translator:uav_address
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                        // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> Green_LEDs_avalon_parallel_port_slave_translator:uav_write
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                         // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Green_LEDs_avalon_parallel_port_slave_translator:uav_lock
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                         // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> Green_LEDs_avalon_parallel_port_slave_translator:uav_read
	wire   [31:0] green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                     // Green_LEDs_avalon_parallel_port_slave_translator:uav_readdata -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                // Green_LEDs_avalon_parallel_port_slave_translator:uav_readdatavalid -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                  // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Green_LEDs_avalon_parallel_port_slave_translator:uav_debugaccess
	wire    [3:0] green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                   // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Green_LEDs_avalon_parallel_port_slave_translator:uav_byteenable
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;           // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                 // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;         // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                  // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                 // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;        // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;              // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;      // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;               // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;              // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;            // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;             // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;            // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // HEX3_HEX0_avalon_parallel_port_slave_translator:uav_waitrequest -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> HEX3_HEX0_avalon_parallel_port_slave_translator:uav_burstcount
	wire   [31:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                     // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> HEX3_HEX0_avalon_parallel_port_slave_translator:uav_writedata
	wire   [28:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                       // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> HEX3_HEX0_avalon_parallel_port_slave_translator:uav_address
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                         // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> HEX3_HEX0_avalon_parallel_port_slave_translator:uav_write
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                          // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> HEX3_HEX0_avalon_parallel_port_slave_translator:uav_lock
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                          // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> HEX3_HEX0_avalon_parallel_port_slave_translator:uav_read
	wire   [31:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                      // HEX3_HEX0_avalon_parallel_port_slave_translator:uav_readdata -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // HEX3_HEX0_avalon_parallel_port_slave_translator:uav_readdatavalid -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> HEX3_HEX0_avalon_parallel_port_slave_translator:uav_debugaccess
	wire    [3:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> HEX3_HEX0_avalon_parallel_port_slave_translator:uav_byteenable
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                   // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Slider_switches_avalon_parallel_port_slave_translator:uav_waitrequest -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Slider_switches_avalon_parallel_port_slave_translator:uav_burstcount
	wire   [31:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Slider_switches_avalon_parallel_port_slave_translator:uav_writedata
	wire   [28:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> Slider_switches_avalon_parallel_port_slave_translator:uav_address
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> Slider_switches_avalon_parallel_port_slave_translator:uav_write
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Slider_switches_avalon_parallel_port_slave_translator:uav_lock
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> Slider_switches_avalon_parallel_port_slave_translator:uav_read
	wire   [31:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // Slider_switches_avalon_parallel_port_slave_translator:uav_readdata -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Slider_switches_avalon_parallel_port_slave_translator:uav_readdatavalid -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Slider_switches_avalon_parallel_port_slave_translator:uav_debugaccess
	wire    [3:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Slider_switches_avalon_parallel_port_slave_translator:uav_byteenable
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // Pushbuttons_avalon_parallel_port_slave_translator:uav_waitrequest -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Pushbuttons_avalon_parallel_port_slave_translator:uav_burstcount
	wire   [31:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                   // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Pushbuttons_avalon_parallel_port_slave_translator:uav_writedata
	wire   [28:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                     // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> Pushbuttons_avalon_parallel_port_slave_translator:uav_address
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                       // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> Pushbuttons_avalon_parallel_port_slave_translator:uav_write
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                        // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Pushbuttons_avalon_parallel_port_slave_translator:uav_lock
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                        // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> Pushbuttons_avalon_parallel_port_slave_translator:uav_read
	wire   [31:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                    // Pushbuttons_avalon_parallel_port_slave_translator:uav_readdata -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // Pushbuttons_avalon_parallel_port_slave_translator:uav_readdatavalid -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Pushbuttons_avalon_parallel_port_slave_translator:uav_debugaccess
	wire    [3:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Pushbuttons_avalon_parallel_port_slave_translator:uav_byteenable
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                 // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;               // Expansion_JP1_avalon_parallel_port_slave_translator:uav_waitrequest -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Expansion_JP1_avalon_parallel_port_slave_translator:uav_burstcount
	wire   [31:0] expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                 // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Expansion_JP1_avalon_parallel_port_slave_translator:uav_writedata
	wire   [28:0] expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                   // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> Expansion_JP1_avalon_parallel_port_slave_translator:uav_address
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                     // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> Expansion_JP1_avalon_parallel_port_slave_translator:uav_write
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                      // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Expansion_JP1_avalon_parallel_port_slave_translator:uav_lock
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                      // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> Expansion_JP1_avalon_parallel_port_slave_translator:uav_read
	wire   [31:0] expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                  // Expansion_JP1_avalon_parallel_port_slave_translator:uav_readdata -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;             // Expansion_JP1_avalon_parallel_port_slave_translator:uav_readdatavalid -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;               // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Expansion_JP1_avalon_parallel_port_slave_translator:uav_debugaccess
	wire    [3:0] expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Expansion_JP1_avalon_parallel_port_slave_translator:uav_byteenable
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;        // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;              // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;      // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;               // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;              // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;     // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;           // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;   // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;            // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;           // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;         // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;          // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;         // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;               // Expansion_JP2_avalon_parallel_port_slave_translator:uav_waitrequest -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Expansion_JP2_avalon_parallel_port_slave_translator:uav_burstcount
	wire   [31:0] expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                 // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Expansion_JP2_avalon_parallel_port_slave_translator:uav_writedata
	wire   [28:0] expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                   // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> Expansion_JP2_avalon_parallel_port_slave_translator:uav_address
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                     // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> Expansion_JP2_avalon_parallel_port_slave_translator:uav_write
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                      // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Expansion_JP2_avalon_parallel_port_slave_translator:uav_lock
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                      // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> Expansion_JP2_avalon_parallel_port_slave_translator:uav_read
	wire   [31:0] expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                  // Expansion_JP2_avalon_parallel_port_slave_translator:uav_readdata -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;             // Expansion_JP2_avalon_parallel_port_slave_translator:uav_readdatavalid -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;               // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Expansion_JP2_avalon_parallel_port_slave_translator:uav_debugaccess
	wire    [3:0] expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Expansion_JP2_avalon_parallel_port_slave_translator:uav_byteenable
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;        // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;              // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;      // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;               // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;              // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;     // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;           // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;   // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;            // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;           // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;         // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;          // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;         // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // Serial_port_avalon_rs232_slave_translator:uav_waitrequest -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Serial_port_avalon_rs232_slave_translator:uav_burstcount
	wire   [31:0] serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                           // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Serial_port_avalon_rs232_slave_translator:uav_writedata
	wire   [28:0] serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_address;                             // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_address -> Serial_port_avalon_rs232_slave_translator:uav_address
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_write;                               // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_write -> Serial_port_avalon_rs232_slave_translator:uav_write
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Serial_port_avalon_rs232_slave_translator:uav_lock
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_read;                                // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_read -> Serial_port_avalon_rs232_slave_translator:uav_read
	wire   [31:0] serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                            // Serial_port_avalon_rs232_slave_translator:uav_readdata -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // Serial_port_avalon_rs232_slave_translator:uav_readdatavalid -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Serial_port_avalon_rs232_slave_translator:uav_debugaccess
	wire    [3:0] serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Serial_port_avalon_rs232_slave_translator:uav_byteenable
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                         // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // Onchip_memory_SRAM_s2_translator:uav_waitrequest -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:m0_burstcount -> Onchip_memory_SRAM_s2_translator:uav_burstcount
	wire   [31:0] onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:m0_writedata -> Onchip_memory_SRAM_s2_translator:uav_writedata
	wire   [28:0] onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_address;                                      // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:m0_address -> Onchip_memory_SRAM_s2_translator:uav_address
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_write;                                        // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:m0_write -> Onchip_memory_SRAM_s2_translator:uav_write
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_lock;                                         // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:m0_lock -> Onchip_memory_SRAM_s2_translator:uav_lock
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_read;                                         // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:m0_read -> Onchip_memory_SRAM_s2_translator:uav_read
	wire   [31:0] onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // Onchip_memory_SRAM_s2_translator:uav_readdata -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // Onchip_memory_SRAM_s2_translator:uav_readdatavalid -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Onchip_memory_SRAM_s2_translator:uav_debugaccess
	wire    [3:0] onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:m0_byteenable -> Onchip_memory_SRAM_s2_translator:uav_byteenable
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rf_source_valid -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rf_source_data -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                                      // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                              // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [103:0] cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                                       // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                                      // addr_router:sink_ready -> cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                       // cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                             // cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                                     // cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [103:0] cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                                              // cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                             // addr_router_001:sink_ready -> cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                                        // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [103:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router:sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                       // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                             // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                     // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [103:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data;                                              // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                             // id_router_001:sink_ready -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                               // sdram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                     // sdram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                             // sdram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire   [85:0] sdram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                      // sdram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                     // id_router_002:sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [103:0] onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_003:sink_ready -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                       // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_rp_valid;                                             // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                     // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [103:0] onchip_memory_s2_translator_avalon_universal_slave_0_agent_rp_data;                                              // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          onchip_memory_s2_translator_avalon_universal_slave_0_agent_rp_ready;                                             // id_router_004:sink_ready -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                  // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [103:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                                   // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_005:sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // Interval_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                            // Interval_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // Interval_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [103:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                             // Interval_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_006:sink_ready -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [103:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_007:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                  // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                        // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [103:0] green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                         // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                        // id_router_008:sink_ready -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                         // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [103:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                          // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_009:sink_ready -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [103:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_010:sink_ready -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                       // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [103:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                        // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router_011:sink_ready -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;               // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                     // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;             // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [103:0] expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                      // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                     // id_router_012:sink_ready -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;               // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                     // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;             // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [103:0] expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                      // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                     // id_router_013:sink_ready -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_valid;                               // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [103:0] serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_data;                                // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_014:sink_ready -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rp_valid;                                        // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [103:0] onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rp_data;                                         // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_015:sink_ready -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:rp_ready
	wire          burst_adapter_source0_endofpacket;                                                                               // burst_adapter:source0_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                                     // burst_adapter:source0_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                             // burst_adapter:source0_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [85:0] burst_adapter_source0_data;                                                                                      // burst_adapter:source0_data -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                                     // sdram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [15:0] burst_adapter_source0_channel;                                                                                   // burst_adapter:source0_channel -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                                  // rst_controller:reset_out -> [Expansion_JP1:reset, Expansion_JP1_avalon_parallel_port_slave_translator:reset, Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Expansion_JP2:reset, Expansion_JP2_avalon_parallel_port_slave_translator:reset, Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Green_LEDs:reset, Green_LEDs_avalon_parallel_port_slave_translator:reset, Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, HEX3_HEX0:reset, HEX3_HEX0_avalon_parallel_port_slave_translator:reset, HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Interval_timer:reset_n, Interval_timer_s1_translator:reset, Interval_timer_s1_translator_avalon_universal_slave_0_agent:reset, Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, JTAG_UART:rst_n, JTAG_UART_avalon_jtag_slave_translator:reset, JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Onchip_memory:reset, Onchip_memory:reset2, Onchip_memory_SRAM:reset, Onchip_memory_SRAM:reset2, Onchip_memory_SRAM_s1_translator:reset, Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:reset, Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Onchip_memory_SRAM_s2_translator:reset, Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:reset, Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Onchip_memory_s1_translator:reset, Onchip_memory_s1_translator_avalon_universal_slave_0_agent:reset, Onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Onchip_memory_s2_translator:reset, Onchip_memory_s2_translator_avalon_universal_slave_0_agent:reset, Onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Pushbuttons:reset, Pushbuttons_avalon_parallel_port_slave_translator:reset, Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Serial_port:reset, Serial_port_avalon_rs232_slave_translator:reset, Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:reset, Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Slider_switches:reset, Slider_switches_avalon_parallel_port_slave_translator:reset, Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, burst_adapter:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_002:reset, cpu:reset_n, cpu_data_master_translator:reset, cpu_data_master_translator_avalon_universal_master_0_agent:reset, cpu_instruction_master_translator:reset, cpu_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_jtag_debug_module_translator:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, irq_mapper:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sdram:reset_n, sdram_s1_translator:reset, sdram_s1_translator_avalon_universal_slave_0_agent:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid:reset_n, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset]
	wire          cpu_jtag_debug_module_reset_reset;                                                                               // cpu:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire          cmd_xbar_demux_src0_endofpacket;                                                                                 // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                                       // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                               // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [103:0] cmd_xbar_demux_src0_data;                                                                                        // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [15:0] cmd_xbar_demux_src0_channel;                                                                                     // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                                       // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                                 // cmd_xbar_demux:src1_endofpacket -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                                       // cmd_xbar_demux:src1_valid -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                               // cmd_xbar_demux:src1_startofpacket -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_src1_data;                                                                                        // cmd_xbar_demux:src1_data -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_src1_channel;                                                                                     // cmd_xbar_demux:src1_channel -> Onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_src2_endofpacket;                                                                                 // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                                       // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                               // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [103:0] cmd_xbar_demux_src2_data;                                                                                        // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire   [15:0] cmd_xbar_demux_src2_channel;                                                                                     // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_src2_ready;                                                                                       // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire          cmd_xbar_demux_src3_endofpacket;                                                                                 // cmd_xbar_demux:src3_endofpacket -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                                       // cmd_xbar_demux:src3_valid -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                                               // cmd_xbar_demux:src3_startofpacket -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_src3_data;                                                                                        // cmd_xbar_demux:src3_data -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_src3_channel;                                                                                     // cmd_xbar_demux:src3_channel -> Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                             // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                                   // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                           // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src0_data;                                                                                    // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [15:0] cmd_xbar_demux_001_src0_channel;                                                                                 // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                                   // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                             // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                                   // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_002:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                           // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src1_data;                                                                                    // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_002:sink1_data
	wire   [15:0] cmd_xbar_demux_001_src1_channel;                                                                                 // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                                   // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                             // cmd_xbar_demux_001:src2_endofpacket -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                                   // cmd_xbar_demux_001:src2_valid -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                           // cmd_xbar_demux_001:src2_startofpacket -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src2_data;                                                                                    // cmd_xbar_demux_001:src2_data -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src2_channel;                                                                                 // cmd_xbar_demux_001:src2_channel -> Onchip_memory_s2_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                             // cmd_xbar_demux_001:src3_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                                   // cmd_xbar_demux_001:src3_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                                           // cmd_xbar_demux_001:src3_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src3_data;                                                                                    // cmd_xbar_demux_001:src3_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src3_channel;                                                                                 // cmd_xbar_demux_001:src3_channel -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                             // cmd_xbar_demux_001:src4_endofpacket -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                                   // cmd_xbar_demux_001:src4_valid -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                                           // cmd_xbar_demux_001:src4_startofpacket -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src4_data;                                                                                    // cmd_xbar_demux_001:src4_data -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src4_channel;                                                                                 // cmd_xbar_demux_001:src4_channel -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                             // cmd_xbar_demux_001:src5_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                                   // cmd_xbar_demux_001:src5_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                                           // cmd_xbar_demux_001:src5_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src5_data;                                                                                    // cmd_xbar_demux_001:src5_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src5_channel;                                                                                 // cmd_xbar_demux_001:src5_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                                             // cmd_xbar_demux_001:src6_endofpacket -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                                   // cmd_xbar_demux_001:src6_valid -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                                           // cmd_xbar_demux_001:src6_startofpacket -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src6_data;                                                                                    // cmd_xbar_demux_001:src6_data -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src6_channel;                                                                                 // cmd_xbar_demux_001:src6_channel -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                                             // cmd_xbar_demux_001:src7_endofpacket -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                                   // cmd_xbar_demux_001:src7_valid -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                                           // cmd_xbar_demux_001:src7_startofpacket -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src7_data;                                                                                    // cmd_xbar_demux_001:src7_data -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src7_channel;                                                                                 // cmd_xbar_demux_001:src7_channel -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src8_endofpacket;                                                                             // cmd_xbar_demux_001:src8_endofpacket -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src8_valid;                                                                                   // cmd_xbar_demux_001:src8_valid -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src8_startofpacket;                                                                           // cmd_xbar_demux_001:src8_startofpacket -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src8_data;                                                                                    // cmd_xbar_demux_001:src8_data -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src8_channel;                                                                                 // cmd_xbar_demux_001:src8_channel -> Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src9_endofpacket;                                                                             // cmd_xbar_demux_001:src9_endofpacket -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src9_valid;                                                                                   // cmd_xbar_demux_001:src9_valid -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src9_startofpacket;                                                                           // cmd_xbar_demux_001:src9_startofpacket -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src9_data;                                                                                    // cmd_xbar_demux_001:src9_data -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src9_channel;                                                                                 // cmd_xbar_demux_001:src9_channel -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src10_endofpacket;                                                                            // cmd_xbar_demux_001:src10_endofpacket -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src10_valid;                                                                                  // cmd_xbar_demux_001:src10_valid -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src10_startofpacket;                                                                          // cmd_xbar_demux_001:src10_startofpacket -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src10_data;                                                                                   // cmd_xbar_demux_001:src10_data -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src10_channel;                                                                                // cmd_xbar_demux_001:src10_channel -> Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src11_endofpacket;                                                                            // cmd_xbar_demux_001:src11_endofpacket -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src11_valid;                                                                                  // cmd_xbar_demux_001:src11_valid -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src11_startofpacket;                                                                          // cmd_xbar_demux_001:src11_startofpacket -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src11_data;                                                                                   // cmd_xbar_demux_001:src11_data -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src11_channel;                                                                                // cmd_xbar_demux_001:src11_channel -> Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src12_endofpacket;                                                                            // cmd_xbar_demux_001:src12_endofpacket -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src12_valid;                                                                                  // cmd_xbar_demux_001:src12_valid -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src12_startofpacket;                                                                          // cmd_xbar_demux_001:src12_startofpacket -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src12_data;                                                                                   // cmd_xbar_demux_001:src12_data -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src12_channel;                                                                                // cmd_xbar_demux_001:src12_channel -> Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src13_endofpacket;                                                                            // cmd_xbar_demux_001:src13_endofpacket -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src13_valid;                                                                                  // cmd_xbar_demux_001:src13_valid -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src13_startofpacket;                                                                          // cmd_xbar_demux_001:src13_startofpacket -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src13_data;                                                                                   // cmd_xbar_demux_001:src13_data -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src13_channel;                                                                                // cmd_xbar_demux_001:src13_channel -> Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                                                 // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                                       // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                               // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [103:0] rsp_xbar_demux_src0_data;                                                                                        // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [15:0] rsp_xbar_demux_src0_channel;                                                                                     // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                                       // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                                 // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                                       // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                               // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [103:0] rsp_xbar_demux_src1_data;                                                                                        // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [15:0] rsp_xbar_demux_src1_channel;                                                                                     // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                                       // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                             // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                                   // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                           // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [103:0] rsp_xbar_demux_001_src0_data;                                                                                    // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [15:0] rsp_xbar_demux_001_src0_channel;                                                                                 // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                                   // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                             // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                                   // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                           // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [103:0] rsp_xbar_demux_002_src0_data;                                                                                    // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [15:0] rsp_xbar_demux_002_src0_channel;                                                                                 // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                                   // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                                             // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                                   // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                                           // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [103:0] rsp_xbar_demux_002_src1_data;                                                                                    // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [15:0] rsp_xbar_demux_002_src1_channel;                                                                                 // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                                   // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_002:src1_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                             // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                                   // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                           // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [103:0] rsp_xbar_demux_003_src0_data;                                                                                    // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire   [15:0] rsp_xbar_demux_003_src0_channel;                                                                                 // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                                   // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                             // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                                   // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                           // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [103:0] rsp_xbar_demux_004_src0_data;                                                                                    // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink2_data
	wire   [15:0] rsp_xbar_demux_004_src0_channel;                                                                                 // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                                   // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                             // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                                   // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                           // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [103:0] rsp_xbar_demux_005_src0_data;                                                                                    // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink3_data
	wire   [15:0] rsp_xbar_demux_005_src0_channel;                                                                                 // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                                   // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                             // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                                   // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                           // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [103:0] rsp_xbar_demux_006_src0_data;                                                                                    // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink4_data
	wire   [15:0] rsp_xbar_demux_006_src0_channel;                                                                                 // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                                   // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                             // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                                   // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                           // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [103:0] rsp_xbar_demux_007_src0_data;                                                                                    // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink5_data
	wire   [15:0] rsp_xbar_demux_007_src0_channel;                                                                                 // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                                   // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                             // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                                   // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                           // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [103:0] rsp_xbar_demux_008_src0_data;                                                                                    // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink6_data
	wire   [15:0] rsp_xbar_demux_008_src0_channel;                                                                                 // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                                   // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                             // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                                   // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                           // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [103:0] rsp_xbar_demux_009_src0_data;                                                                                    // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink7_data
	wire   [15:0] rsp_xbar_demux_009_src0_channel;                                                                                 // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                                   // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                             // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                                   // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                           // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [103:0] rsp_xbar_demux_010_src0_data;                                                                                    // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink8_data
	wire   [15:0] rsp_xbar_demux_010_src0_channel;                                                                                 // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                                   // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                             // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                                   // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                           // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [103:0] rsp_xbar_demux_011_src0_data;                                                                                    // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink9_data
	wire   [15:0] rsp_xbar_demux_011_src0_channel;                                                                                 // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                                   // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                             // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                                   // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                                           // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [103:0] rsp_xbar_demux_012_src0_data;                                                                                    // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink10_data
	wire   [15:0] rsp_xbar_demux_012_src0_channel;                                                                                 // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                                   // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                             // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                                   // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                                           // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [103:0] rsp_xbar_demux_013_src0_data;                                                                                    // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_001:sink11_data
	wire   [15:0] rsp_xbar_demux_013_src0_channel;                                                                                 // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                                   // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_013:src0_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                                             // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                                   // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_001:sink12_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                                           // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [103:0] rsp_xbar_demux_014_src0_data;                                                                                    // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_001:sink12_data
	wire   [15:0] rsp_xbar_demux_014_src0_channel;                                                                                 // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_001:sink12_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                                   // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                                             // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                                   // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_001:sink13_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                                           // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [103:0] rsp_xbar_demux_015_src0_data;                                                                                    // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_001:sink13_data
	wire   [15:0] rsp_xbar_demux_015_src0_channel;                                                                                 // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_001:sink13_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                                   // rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_015:src0_ready
	wire          addr_router_src_endofpacket;                                                                                     // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                                                           // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                                                   // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [103:0] addr_router_src_data;                                                                                            // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [15:0] addr_router_src_channel;                                                                                         // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                                                           // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                                    // rsp_xbar_mux:src_endofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                          // rsp_xbar_mux:src_valid -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                                  // rsp_xbar_mux:src_startofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [103:0] rsp_xbar_mux_src_data;                                                                                           // rsp_xbar_mux:src_data -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] rsp_xbar_mux_src_channel;                                                                                        // rsp_xbar_mux:src_channel -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_src_ready;                                                                                          // cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                                 // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                                       // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                               // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [103:0] addr_router_001_src_data;                                                                                        // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [15:0] addr_router_001_src_channel;                                                                                     // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                                       // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                                // rsp_xbar_mux_001:src_endofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                                      // rsp_xbar_mux_001:src_valid -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                              // rsp_xbar_mux_001:src_startofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [103:0] rsp_xbar_mux_001_src_data;                                                                                       // rsp_xbar_mux_001:src_data -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] rsp_xbar_mux_001_src_channel;                                                                                    // rsp_xbar_mux_001:src_channel -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                                      // cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                                    // cmd_xbar_mux:src_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                          // cmd_xbar_mux:src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                                  // cmd_xbar_mux:src_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_mux_src_data;                                                                                           // cmd_xbar_mux:src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_mux_src_channel;                                                                                        // cmd_xbar_mux:src_channel -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                                       // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                             // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                                     // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [103:0] id_router_src_data;                                                                                              // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [15:0] id_router_src_channel;                                                                                           // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                             // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_demux_src1_ready;                                                                                       // Onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src1_ready
	wire          id_router_001_src_endofpacket;                                                                                   // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                                         // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                                 // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [103:0] id_router_001_src_data;                                                                                          // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [15:0] id_router_001_src_channel;                                                                                       // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                                         // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_demux_src3_ready;                                                                                       // Onchip_memory_SRAM_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src3_ready
	wire          id_router_003_src_endofpacket;                                                                                   // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                         // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                                 // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [103:0] id_router_003_src_data;                                                                                          // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [15:0] id_router_003_src_channel;                                                                                       // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                         // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_001_src2_ready;                                                                                   // Onchip_memory_s2_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src2_ready
	wire          id_router_004_src_endofpacket;                                                                                   // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                         // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                                 // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [103:0] id_router_004_src_data;                                                                                          // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [15:0] id_router_004_src_channel;                                                                                       // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                         // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_demux_001_src3_ready;                                                                                   // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire          id_router_005_src_endofpacket;                                                                                   // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                                         // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                                 // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [103:0] id_router_005_src_data;                                                                                          // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [15:0] id_router_005_src_channel;                                                                                       // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                                         // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_001_src4_ready;                                                                                   // Interval_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire          id_router_006_src_endofpacket;                                                                                   // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                         // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                                 // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [103:0] id_router_006_src_data;                                                                                          // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [15:0] id_router_006_src_channel;                                                                                       // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                         // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_001_src5_ready;                                                                                   // sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire          id_router_007_src_endofpacket;                                                                                   // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                         // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                                 // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [103:0] id_router_007_src_data;                                                                                          // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [15:0] id_router_007_src_channel;                                                                                       // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                         // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_001_src6_ready;                                                                                   // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire          id_router_008_src_endofpacket;                                                                                   // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                         // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                                 // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [103:0] id_router_008_src_data;                                                                                          // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [15:0] id_router_008_src_channel;                                                                                       // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                         // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_demux_001_src7_ready;                                                                                   // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire          id_router_009_src_endofpacket;                                                                                   // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                         // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                                 // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [103:0] id_router_009_src_data;                                                                                          // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [15:0] id_router_009_src_channel;                                                                                       // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                         // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_001_src8_ready;                                                                                   // Slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire          id_router_010_src_endofpacket;                                                                                   // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                                         // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                                 // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [103:0] id_router_010_src_data;                                                                                          // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [15:0] id_router_010_src_channel;                                                                                       // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                                         // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_001_src9_ready;                                                                                   // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	wire          id_router_011_src_endofpacket;                                                                                   // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                                         // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                                 // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [103:0] id_router_011_src_data;                                                                                          // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [15:0] id_router_011_src_channel;                                                                                       // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                                         // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_demux_001_src10_ready;                                                                                  // Expansion_JP1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	wire          id_router_012_src_endofpacket;                                                                                   // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                                         // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                                 // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [103:0] id_router_012_src_data;                                                                                          // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [15:0] id_router_012_src_channel;                                                                                       // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                                         // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          cmd_xbar_demux_001_src11_ready;                                                                                  // Expansion_JP2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	wire          id_router_013_src_endofpacket;                                                                                   // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                                         // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                                 // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [103:0] id_router_013_src_data;                                                                                          // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [15:0] id_router_013_src_channel;                                                                                       // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                                         // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_demux_001_src12_ready;                                                                                  // Serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	wire          id_router_014_src_endofpacket;                                                                                   // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                                         // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                                 // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [103:0] id_router_014_src_data;                                                                                          // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [15:0] id_router_014_src_channel;                                                                                       // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                                         // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          cmd_xbar_demux_001_src13_ready;                                                                                  // Onchip_memory_SRAM_s2_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src13_ready
	wire          id_router_015_src_endofpacket;                                                                                   // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                                         // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                                 // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [103:0] id_router_015_src_data;                                                                                          // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [15:0] id_router_015_src_channel;                                                                                       // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                                         // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                                // cmd_xbar_mux_002:src_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                                      // cmd_xbar_mux_002:src_valid -> width_adapter:in_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                                              // cmd_xbar_mux_002:src_startofpacket -> width_adapter:in_startofpacket
	wire  [103:0] cmd_xbar_mux_002_src_data;                                                                                       // cmd_xbar_mux_002:src_data -> width_adapter:in_data
	wire   [15:0] cmd_xbar_mux_002_src_channel;                                                                                    // cmd_xbar_mux_002:src_channel -> width_adapter:in_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                                      // width_adapter:in_ready -> cmd_xbar_mux_002:src_ready
	wire          width_adapter_src_endofpacket;                                                                                   // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                                         // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                                 // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [85:0] width_adapter_src_data;                                                                                          // width_adapter:out_data -> burst_adapter:sink0_data
	wire          width_adapter_src_ready;                                                                                         // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire   [15:0] width_adapter_src_channel;                                                                                       // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire          id_router_002_src_endofpacket;                                                                                   // id_router_002:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_002_src_valid;                                                                                         // id_router_002:src_valid -> width_adapter_001:in_valid
	wire          id_router_002_src_startofpacket;                                                                                 // id_router_002:src_startofpacket -> width_adapter_001:in_startofpacket
	wire   [85:0] id_router_002_src_data;                                                                                          // id_router_002:src_data -> width_adapter_001:in_data
	wire   [15:0] id_router_002_src_channel;                                                                                       // id_router_002:src_channel -> width_adapter_001:in_channel
	wire          id_router_002_src_ready;                                                                                         // width_adapter_001:in_ready -> id_router_002:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                               // width_adapter_001:out_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                                     // width_adapter_001:out_valid -> rsp_xbar_demux_002:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                                             // width_adapter_001:out_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [103:0] width_adapter_001_src_data;                                                                                      // width_adapter_001:out_data -> rsp_xbar_demux_002:sink_data
	wire          width_adapter_001_src_ready;                                                                                     // rsp_xbar_demux_002:sink_ready -> width_adapter_001:out_ready
	wire   [15:0] width_adapter_001_src_channel;                                                                                   // width_adapter_001:out_channel -> rsp_xbar_demux_002:sink_channel
	wire          irq_mapper_receiver0_irq;                                                                                        // JTAG_UART:av_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                                        // Interval_timer:irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                                                        // Serial_port:irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                                                        // Pushbuttons:irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                                                                        // Expansion_JP1:irq -> irq_mapper:receiver4_irq
	wire          irq_mapper_receiver5_irq;                                                                                        // Expansion_JP2:irq -> irq_mapper:receiver5_irq
	wire   [31:0] cpu_d_irq_irq;                                                                                                   // irq_mapper:sender_irq -> cpu:d_irq

	nios_system_Onchip_memory onchip_memory (
		.clk         (clk),                                                        //   clk1.clk
		.address     (onchip_memory_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken       (onchip_memory_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect  (onchip_memory_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write       (onchip_memory_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata    (onchip_memory_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata   (onchip_memory_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable  (onchip_memory_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                             // reset1.reset
		.address2    (onchip_memory_s2_translator_avalon_anti_slave_0_address),    //     s2.address
		.chipselect2 (onchip_memory_s2_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken2      (onchip_memory_s2_translator_avalon_anti_slave_0_clken),      //       .clken
		.write2      (onchip_memory_s2_translator_avalon_anti_slave_0_write),      //       .write
		.readdata2   (onchip_memory_s2_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata2  (onchip_memory_s2_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable2 (onchip_memory_s2_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.clk2        (clk),                                                        //   clk2.clk
		.reset2      (rst_controller_reset_out_reset)                              // reset2.reset
	);

	nios_system_JTAG_UART jtag_uart (
		.clk            (clk),                                                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                //               irq.irq
	);

	nios_system_Interval_timer interval_timer (
		.clk        (clk),                                                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                             // reset.reset_n
		.address    (interval_timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (interval_timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (interval_timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (interval_timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~interval_timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                                     //   irq.irq
	);

	nios_system_sdram sdram (
		.clk            (clk),                                                   //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                       // reset.reset_n
		.az_addr        (sdram_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (zs_addr_from_the_sdram),                                //  wire.export
		.zs_ba          (zs_ba_from_the_sdram),                                  //      .export
		.zs_cas_n       (zs_cas_n_from_the_sdram),                               //      .export
		.zs_cke         (zs_cke_from_the_sdram),                                 //      .export
		.zs_cs_n        (zs_cs_n_from_the_sdram),                                //      .export
		.zs_dq          (zs_dq_to_and_from_the_sdram),                           //      .export
		.zs_dqm         (zs_dqm_from_the_sdram),                                 //      .export
		.zs_ras_n       (zs_ras_n_from_the_sdram),                               //      .export
		.zs_we_n        (zs_we_n_from_the_sdram)                                 //      .export
	);

	nios_system_Green_LEDs green_leds (
		.clk        (clk),                                                                             //                clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                                  //          clock_reset_reset.reset
		.address    (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.LEDG       (LEDG_from_the_Green_LEDs)                                                         //         external_interface.export
	);

	nios_system_HEX3_HEX0 hex3_hex0 (
		.clk        (clk),                                                                            //                clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                                 //          clock_reset_reset.reset
		.address    (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.HEX0       (HEX0_from_the_HEX3_HEX0),                                                        //         external_interface.export
		.HEX1       (HEX1_from_the_HEX3_HEX0),                                                        //                           .export
		.HEX2       (HEX2_from_the_HEX3_HEX0),                                                        //                           .export
		.HEX3       (HEX3_from_the_HEX3_HEX0)                                                         //                           .export
	);

	nios_system_Slider_switches slider_switches (
		.clk        (clk),                                                                                  //                clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                                       //          clock_reset_reset.reset
		.address    (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.SW         (SW_to_the_Slider_switches)                                                             //         external_interface.export
	);

	nios_system_Pushbuttons pushbuttons (
		.clk        (clk),                                                                              //                clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                                   //          clock_reset_reset.reset
		.address    (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.KEY        (KEY_to_the_Pushbuttons),                                                           //         external_interface.export
		.irq        (irq_mapper_receiver3_irq)                                                          //                  interrupt.irq
	);

	nios_system_Expansion_JP1 expansion_jp1 (
		.clk        (clk),                                                                                //                clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                                     //          clock_reset_reset.reset
		.address    (expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.GPIO_0     (GPIO_0_to_and_from_the_Expansion_JP1),                                               //         external_interface.export
		.irq        (irq_mapper_receiver4_irq)                                                            //                  interrupt.irq
	);

	nios_system_Expansion_JP2 expansion_jp2 (
		.clk        (clk),                                                                                //                clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                                     //          clock_reset_reset.reset
		.address    (expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.GPIO_1     (GPIO_1_to_and_from_the_Expansion_JP2),                                               //         external_interface.export
		.irq        (irq_mapper_receiver5_irq)                                                            //                  interrupt.irq
	);

	nios_system_Serial_port serial_port (
		.clk        (clk),                                                                      //        clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                           //  clock_reset_reset.reset
		.address    (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_address),    // avalon_rs232_slave.address
		.chipselect (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.byteenable (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_byteenable), //                   .byteenable
		.read       (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_read),       //                   .read
		.write      (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_write),      //                   .write
		.writedata  (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.readdata   (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver2_irq),                                                 //          interrupt.irq
		.UART_RXD   (UART_RXD_to_the_Serial_port),                                              // external_interface.export
		.UART_TXD   (UART_TXD_from_the_Serial_port)                                             //                   .export
	);

	nios_system_Onchip_memory_SRAM onchip_memory_sram (
		.clk         (clk),                                                             //   clk1.clk
		.address     (onchip_memory_sram_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken       (onchip_memory_sram_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect  (onchip_memory_sram_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write       (onchip_memory_sram_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata    (onchip_memory_sram_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata   (onchip_memory_sram_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable  (onchip_memory_sram_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                                  // reset1.reset
		.address2    (onchip_memory_sram_s2_translator_avalon_anti_slave_0_address),    //     s2.address
		.chipselect2 (onchip_memory_sram_s2_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken2      (onchip_memory_sram_s2_translator_avalon_anti_slave_0_clken),      //       .clken
		.write2      (onchip_memory_sram_s2_translator_avalon_anti_slave_0_write),      //       .write
		.readdata2   (onchip_memory_sram_s2_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata2  (onchip_memory_sram_s2_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable2 (onchip_memory_sram_s2_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.clk2        (clk),                                                             //   clk2.clk
		.reset2      (rst_controller_reset_out_reset)                                   // reset2.reset
	);

	nios_system_cpu cpu (
		.clk                                   (clk),                                                              //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                  //                   reset_n.reset_n
		.d_address                             (cpu_data_master_address),                                          //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (cpu_data_master_read),                                             //                          .read
		.d_readdata                            (cpu_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (cpu_data_master_write),                                            //                          .write
		.d_writedata                           (cpu_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                                      //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                               //                          .waitrequest
		.d_irq                                 (cpu_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (cpu_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                  // custom_instruction_master.readra
	);

	nios_system_sysid sysid (
		.clock    (clk),                                                         //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                             //         reset.reset_n
		.readdata (sysid_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (29),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_instruction_master_translator (
		.clk                      (clk),                                                                       //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                            //                     reset.reset
		.uav_address              (cpu_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (cpu_instruction_master_read),                                               //                          .read
		.av_readdata              (cpu_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                      //               (terminated)
		.av_byteenable            (4'b1111),                                                                   //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                      //               (terminated)
		.av_begintransfer         (1'b0),                                                                      //               (terminated)
		.av_chipselect            (1'b0),                                                                      //               (terminated)
		.av_readdatavalid         (),                                                                          //               (terminated)
		.av_write                 (1'b0),                                                                      //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                      //               (terminated)
		.av_lock                  (1'b0),                                                                      //               (terminated)
		.av_debugaccess           (1'b0),                                                                      //               (terminated)
		.uav_clken                (),                                                                          //               (terminated)
		.av_clken                 (1'b1),                                                                      //               (terminated)
		.uav_response             (2'b00),                                                                     //               (terminated)
		.av_response              (),                                                                          //               (terminated)
		.uav_writeresponserequest (),                                                                          //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                      //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                      //               (terminated)
		.av_writeresponsevalid    ()                                                                           //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (29),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (29),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) cpu_data_master_translator (
		.clk                      (clk),                                                                //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                     reset.reset
		.uav_address              (cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (cpu_data_master_read),                                               //                          .read
		.av_readdata              (cpu_data_master_readdata),                                           //                          .readdata
		.av_write                 (cpu_data_master_write),                                              //                          .write
		.av_writedata             (cpu_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                               //               (terminated)
		.av_begintransfer         (1'b0),                                                               //               (terminated)
		.av_chipselect            (1'b0),                                                               //               (terminated)
		.av_readdatavalid         (),                                                                   //               (terminated)
		.av_lock                  (1'b0),                                                               //               (terminated)
		.uav_clken                (),                                                                   //               (terminated)
		.av_clken                 (1'b1),                                                               //               (terminated)
		.uav_response             (2'b00),                                                              //               (terminated)
		.av_response              (),                                                                   //               (terminated)
		.uav_writeresponserequest (),                                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                                               //               (terminated)
		.av_writeresponsevalid    ()                                                                    //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (29),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_jtag_debug_module_translator (
		.clk                      (clk),                                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                   //                    reset.reset
		.uav_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (cpu_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                                 //              (terminated)
		.av_burstcount            (),                                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                                             //              (terminated)
		.av_writebyteenable       (),                                                                                 //              (terminated)
		.av_lock                  (),                                                                                 //              (terminated)
		.av_chipselect            (),                                                                                 //              (terminated)
		.av_clken                 (),                                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                                             //              (terminated)
		.av_outputenable          (),                                                                                 //              (terminated)
		.uav_response             (),                                                                                 //              (terminated)
		.av_response              (2'b00),                                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (11),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (29),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory_s1_translator (
		.clk                      (clk),                                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address              (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_memory_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_memory_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_memory_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_memory_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_memory_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_memory_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_memory_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (29),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_s1_translator (
		.clk                      (clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sdram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sdram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sdram_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sdram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sdram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sdram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (sdram_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (sdram_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (sdram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (11),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (29),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory_sram_s1_translator (
		.clk                      (clk),                                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                   //                    reset.reset
		.uav_address              (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_memory_sram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_memory_sram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_memory_sram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_memory_sram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_memory_sram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_memory_sram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_memory_sram_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                                 //              (terminated)
		.av_begintransfer         (),                                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                                 //              (terminated)
		.av_burstcount            (),                                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                                             //              (terminated)
		.av_waitrequest           (1'b0),                                                                             //              (terminated)
		.av_writebyteenable       (),                                                                                 //              (terminated)
		.av_lock                  (),                                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                                             //              (terminated)
		.av_debugaccess           (),                                                                                 //              (terminated)
		.av_outputenable          (),                                                                                 //              (terminated)
		.uav_response             (),                                                                                 //              (terminated)
		.av_response              (2'b00),                                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (11),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (29),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory_s2_translator (
		.clk                      (clk),                                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address              (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_memory_s2_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_memory_s2_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_memory_s2_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_memory_s2_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_memory_s2_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_memory_s2_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_memory_s2_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (29),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                      (clk),                                                                                    //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_byteenable            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (29),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) interval_timer_s1_translator (
		.clk                      (clk),                                                                          //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                               //                    reset.reset
		.uav_address              (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (interval_timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (interval_timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (interval_timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (interval_timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (interval_timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                             //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (29),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_control_slave_translator (
		.clk                      (clk),                                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sysid_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (sysid_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                               //              (terminated)
		.av_read                  (),                                                                               //              (terminated)
		.av_writedata             (),                                                                               //              (terminated)
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_byteenable            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_chipselect            (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (29),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) green_leds_avalon_parallel_port_slave_translator (
		.clk                      (clk),                                                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                   //                    reset.reset
		.uav_address              (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                                                 //              (terminated)
		.av_burstcount            (),                                                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                             //              (terminated)
		.av_waitrequest           (1'b0),                                                                                             //              (terminated)
		.av_writebyteenable       (),                                                                                                 //              (terminated)
		.av_lock                  (),                                                                                                 //              (terminated)
		.av_clken                 (),                                                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                                                             //              (terminated)
		.av_debugaccess           (),                                                                                                 //              (terminated)
		.av_outputenable          (),                                                                                                 //              (terminated)
		.uav_response             (),                                                                                                 //              (terminated)
		.av_response              (2'b00),                                                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (29),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex3_hex0_avalon_parallel_port_slave_translator (
		.clk                      (clk),                                                                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                  //                    reset.reset
		.uav_address              (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                //              (terminated)
		.av_beginbursttransfer    (),                                                                                                //              (terminated)
		.av_burstcount            (),                                                                                                //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                            //              (terminated)
		.av_waitrequest           (1'b0),                                                                                            //              (terminated)
		.av_writebyteenable       (),                                                                                                //              (terminated)
		.av_lock                  (),                                                                                                //              (terminated)
		.av_clken                 (),                                                                                                //              (terminated)
		.uav_clken                (1'b0),                                                                                            //              (terminated)
		.av_debugaccess           (),                                                                                                //              (terminated)
		.av_outputenable          (),                                                                                                //              (terminated)
		.uav_response             (),                                                                                                //              (terminated)
		.av_response              (2'b00),                                                                                           //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                            //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                //              (terminated)
		.av_writeresponserequest  (),                                                                                                //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (29),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) slider_switches_avalon_parallel_port_slave_translator (
		.clk                      (clk),                                                                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                        //                    reset.reset
		.uav_address              (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                                                      //              (terminated)
		.av_burstcount            (),                                                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                                      //              (terminated)
		.av_lock                  (),                                                                                                      //              (terminated)
		.av_clken                 (),                                                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                                                  //              (terminated)
		.av_debugaccess           (),                                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                                      //              (terminated)
		.uav_response             (),                                                                                                      //              (terminated)
		.av_response              (2'b00),                                                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (29),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pushbuttons_avalon_parallel_port_slave_translator (
		.clk                      (clk),                                                                                               //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                    //                    reset.reset
		.uav_address              (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                                                  //              (terminated)
		.av_burstcount            (),                                                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                                                              //              (terminated)
		.av_writebyteenable       (),                                                                                                  //              (terminated)
		.av_lock                  (),                                                                                                  //              (terminated)
		.av_clken                 (),                                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                                              //              (terminated)
		.av_debugaccess           (),                                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                                  //              (terminated)
		.uav_response             (),                                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (29),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) expansion_jp1_avalon_parallel_port_slave_translator (
		.clk                      (clk),                                                                                                 //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                      //                    reset.reset
		.uav_address              (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (expansion_jp1_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                                    //              (terminated)
		.av_burstcount            (),                                                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                                    //              (terminated)
		.av_lock                  (),                                                                                                    //              (terminated)
		.av_clken                 (),                                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                                //              (terminated)
		.av_debugaccess           (),                                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                                    //              (terminated)
		.uav_response             (),                                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (29),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) expansion_jp2_avalon_parallel_port_slave_translator (
		.clk                      (clk),                                                                                                 //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                      //                    reset.reset
		.uav_address              (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (expansion_jp2_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                                    //              (terminated)
		.av_burstcount            (),                                                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                                    //              (terminated)
		.av_lock                  (),                                                                                                    //              (terminated)
		.av_clken                 (),                                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                                //              (terminated)
		.av_debugaccess           (),                                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                                    //              (terminated)
		.uav_response             (),                                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (29),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) serial_port_avalon_rs232_slave_translator (
		.clk                      (clk),                                                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address              (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                                          //              (terminated)
		.av_burstcount            (),                                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                                          //              (terminated)
		.av_lock                  (),                                                                                          //              (terminated)
		.av_clken                 (),                                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                                      //              (terminated)
		.av_debugaccess           (),                                                                                          //              (terminated)
		.av_outputenable          (),                                                                                          //              (terminated)
		.uav_response             (),                                                                                          //              (terminated)
		.av_response              (2'b00),                                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (11),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (29),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory_sram_s2_translator (
		.clk                      (clk),                                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                   //                    reset.reset
		.uav_address              (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_memory_sram_s2_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_memory_sram_s2_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_memory_sram_s2_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_memory_sram_s2_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_memory_sram_s2_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_memory_sram_s2_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_memory_sram_s2_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                                 //              (terminated)
		.av_begintransfer         (),                                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                                 //              (terminated)
		.av_burstcount            (),                                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                                             //              (terminated)
		.av_waitrequest           (1'b0),                                                                             //              (terminated)
		.av_writebyteenable       (),                                                                                 //              (terminated)
		.av_lock                  (),                                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                                             //              (terminated)
		.av_debugaccess           (),                                                                                 //              (terminated)
		.av_outputenable          (),                                                                                 //              (terminated)
		.uav_response             (),                                                                                 //              (terminated)
		.av_response              (2'b00),                                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                              //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_BEGIN_BURST           (84),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (74),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.PKT_BURST_TYPE_H          (81),
		.PKT_BURST_TYPE_L          (80),
		.PKT_BYTE_CNT_H            (73),
		.PKT_BYTE_CNT_L            (71),
		.PKT_ADDR_H                (64),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (65),
		.PKT_TRANS_POSTED          (66),
		.PKT_TRANS_WRITE           (67),
		.PKT_TRANS_READ            (68),
		.PKT_TRANS_LOCK            (69),
		.PKT_TRANS_EXCLUSIVE       (70),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (90),
		.PKT_THREAD_ID_H           (94),
		.PKT_THREAD_ID_L           (94),
		.PKT_CACHE_H               (101),
		.PKT_CACHE_L               (98),
		.PKT_DATA_SIDEBAND_H       (83),
		.PKT_DATA_SIDEBAND_L       (83),
		.PKT_QOS_H                 (85),
		.PKT_QOS_L                 (85),
		.PKT_ADDR_SIDEBAND_H       (82),
		.PKT_ADDR_SIDEBAND_L       (82),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.ST_DATA_W                 (104),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk),                                                                                //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.av_address              (cpu_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_src_valid),                                                             //        rp.valid
		.rp_data                 (rsp_xbar_mux_src_data),                                                              //          .data
		.rp_channel              (rsp_xbar_mux_src_channel),                                                           //          .channel
		.rp_startofpacket        (rsp_xbar_mux_src_startofpacket),                                                     //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_src_endofpacket),                                                       //          .endofpacket
		.rp_ready                (rsp_xbar_mux_src_ready),                                                             //          .ready
		.av_response             (),                                                                                   // (terminated)
		.av_writeresponserequest (1'b0),                                                                               // (terminated)
		.av_writeresponsevalid   ()                                                                                    // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_BEGIN_BURST           (84),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (74),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.PKT_BURST_TYPE_H          (81),
		.PKT_BURST_TYPE_L          (80),
		.PKT_BYTE_CNT_H            (73),
		.PKT_BYTE_CNT_L            (71),
		.PKT_ADDR_H                (64),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (65),
		.PKT_TRANS_POSTED          (66),
		.PKT_TRANS_WRITE           (67),
		.PKT_TRANS_READ            (68),
		.PKT_TRANS_LOCK            (69),
		.PKT_TRANS_EXCLUSIVE       (70),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (90),
		.PKT_THREAD_ID_H           (94),
		.PKT_THREAD_ID_L           (94),
		.PKT_CACHE_H               (101),
		.PKT_CACHE_L               (98),
		.PKT_DATA_SIDEBAND_H       (83),
		.PKT_DATA_SIDEBAND_L       (83),
		.PKT_QOS_H                 (85),
		.PKT_QOS_L                 (85),
		.PKT_ADDR_SIDEBAND_H       (82),
		.PKT_ADDR_SIDEBAND_L       (82),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.ST_DATA_W                 (104),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk),                                                                         //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.av_address              (cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_001_src_valid),                                                  //        rp.valid
		.rp_data                 (rsp_xbar_mux_001_src_data),                                                   //          .data
		.rp_channel              (rsp_xbar_mux_001_src_channel),                                                //          .channel
		.rp_startofpacket        (rsp_xbar_mux_001_src_startofpacket),                                          //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_001_src_endofpacket),                                            //          .endofpacket
		.rp_ready                (rsp_xbar_mux_001_src_ready),                                                  //          .ready
		.av_response             (),                                                                            // (terminated)
		.av_writeresponserequest (1'b0),                                                                        // (terminated)
		.av_writeresponsevalid   ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (64),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (65),
		.PKT_TRANS_POSTED          (66),
		.PKT_TRANS_WRITE           (67),
		.PKT_TRANS_READ            (68),
		.PKT_TRANS_LOCK            (69),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (74),
		.PKT_BYTE_CNT_H            (73),
		.PKT_BYTE_CNT_L            (71),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                   //                .channel
		.rf_sink_ready           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (64),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (65),
		.PKT_TRANS_POSTED          (66),
		.PKT_TRANS_WRITE           (67),
		.PKT_TRANS_READ            (68),
		.PKT_TRANS_LOCK            (69),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (74),
		.PKT_BYTE_CNT_H            (73),
		.PKT_BYTE_CNT_L            (71),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_memory_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src1_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_src1_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_src1_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_src1_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src1_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src1_channel),                                                           //                .channel
		.rf_sink_ready           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (46),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (47),
		.PKT_TRANS_POSTED          (48),
		.PKT_TRANS_WRITE           (49),
		.PKT_TRANS_READ            (50),
		.PKT_TRANS_LOCK            (51),
		.PKT_SRC_ID_H              (71),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (75),
		.PKT_DEST_ID_L             (72),
		.PKT_BURSTWRAP_H           (58),
		.PKT_BURSTWRAP_L           (56),
		.PKT_BYTE_CNT_H            (55),
		.PKT_BYTE_CNT_L            (53),
		.PKT_PROTECTION_H          (79),
		.PKT_PROTECTION_L          (77),
		.PKT_RESPONSE_STATUS_H     (85),
		.PKT_RESPONSE_STATUS_L     (84),
		.PKT_BURST_SIZE_H          (61),
		.PKT_BURST_SIZE_L          (59),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (86),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                   //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                   //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                    //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                             //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                 //                .channel
		.rf_sink_ready           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (87),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (18),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk),                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                   // (terminated)
		.csr_read          (1'b0),                                                                    // (terminated)
		.csr_write         (1'b0),                                                                    // (terminated)
		.csr_readdata      (),                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                    // (terminated)
		.almost_full_data  (),                                                                        // (terminated)
		.almost_empty_data (),                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                    // (terminated)
		.out_startofpacket (),                                                                        // (terminated)
		.out_endofpacket   (),                                                                        // (terminated)
		.in_empty          (1'b0),                                                                    // (terminated)
		.out_empty         (),                                                                        // (terminated)
		.in_error          (1'b0),                                                                    // (terminated)
		.out_error         (),                                                                        // (terminated)
		.in_channel        (1'b0),                                                                    // (terminated)
		.out_channel       ()                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (64),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (65),
		.PKT_TRANS_POSTED          (66),
		.PKT_TRANS_WRITE           (67),
		.PKT_TRANS_READ            (68),
		.PKT_TRANS_LOCK            (69),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (74),
		.PKT_BYTE_CNT_H            (73),
		.PKT_BYTE_CNT_L            (71),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src3_ready),                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_src3_valid),                                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_src3_data),                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_src3_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src3_endofpacket),                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src3_channel),                                                                //                .channel
		.rf_sink_ready           (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (64),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (65),
		.PKT_TRANS_POSTED          (66),
		.PKT_TRANS_WRITE           (67),
		.PKT_TRANS_READ            (68),
		.PKT_TRANS_LOCK            (69),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (74),
		.PKT_BYTE_CNT_H            (73),
		.PKT_BYTE_CNT_L            (71),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_memory_s2_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory_s2_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src2_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src2_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src2_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src2_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src2_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src2_channel),                                                       //                .channel
		.rf_sink_ready           (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (64),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (65),
		.PKT_TRANS_POSTED          (66),
		.PKT_TRANS_WRITE           (67),
		.PKT_TRANS_READ            (68),
		.PKT_TRANS_LOCK            (69),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (74),
		.PKT_BYTE_CNT_H            (73),
		.PKT_BYTE_CNT_L            (71),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (64),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (65),
		.PKT_TRANS_POSTED          (66),
		.PKT_TRANS_WRITE           (67),
		.PKT_TRANS_READ            (68),
		.PKT_TRANS_LOCK            (69),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (74),
		.PKT_BYTE_CNT_H            (73),
		.PKT_BYTE_CNT_L            (71),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) interval_timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                        //                .channel
		.rf_sink_ready           (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (64),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (65),
		.PKT_TRANS_POSTED          (66),
		.PKT_TRANS_WRITE           (67),
		.PKT_TRANS_READ            (68),
		.PKT_TRANS_LOCK            (69),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (74),
		.PKT_BYTE_CNT_H            (73),
		.PKT_BYTE_CNT_L            (71),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                          //                .channel
		.rf_sink_ready           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (64),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (65),
		.PKT_TRANS_POSTED          (66),
		.PKT_TRANS_WRITE           (67),
		.PKT_TRANS_READ            (68),
		.PKT_TRANS_LOCK            (69),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (74),
		.PKT_BYTE_CNT_H            (73),
		.PKT_BYTE_CNT_L            (71),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                             //       clk_reset.reset
		.m0_address              (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                                            //                .channel
		.rf_sink_ready           (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                             // clk_reset.reset
		.in_data           (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                                       // (terminated)
		.csr_readdata      (),                                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                       // (terminated)
		.almost_full_data  (),                                                                                                           // (terminated)
		.almost_empty_data (),                                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                                       // (terminated)
		.out_empty         (),                                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                                       // (terminated)
		.out_error         (),                                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                                       // (terminated)
		.out_channel       ()                                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (64),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (65),
		.PKT_TRANS_POSTED          (66),
		.PKT_TRANS_WRITE           (67),
		.PKT_TRANS_READ            (68),
		.PKT_TRANS_LOCK            (69),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (74),
		.PKT_BYTE_CNT_H            (73),
		.PKT_BYTE_CNT_L            (71),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                            //       clk_reset.reset
		.m0_address              (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                                           //                .channel
		.rf_sink_ready           (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                     //     (terminated)
		.m0_writeresponserequest (),                                                                                                          //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                       //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                            // clk_reset.reset
		.in_data           (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                                      // (terminated)
		.csr_readdata      (),                                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                      // (terminated)
		.almost_full_data  (),                                                                                                          // (terminated)
		.almost_empty_data (),                                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                                      // (terminated)
		.out_empty         (),                                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                                      // (terminated)
		.out_error         (),                                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                                      // (terminated)
		.out_channel       ()                                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (64),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (65),
		.PKT_TRANS_POSTED          (66),
		.PKT_TRANS_WRITE           (67),
		.PKT_TRANS_READ            (68),
		.PKT_TRANS_LOCK            (69),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (74),
		.PKT_BYTE_CNT_H            (73),
		.PKT_BYTE_CNT_L            (71),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                  //       clk_reset.reset
		.m0_address              (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                                                 //                .channel
		.rf_sink_ready           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                  // clk_reset.reset
		.in_data           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                            // (terminated)
		.almost_full_data  (),                                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                                            // (terminated)
		.out_empty         (),                                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                                            // (terminated)
		.out_error         (),                                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                                            // (terminated)
		.out_channel       ()                                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (64),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (65),
		.PKT_TRANS_POSTED          (66),
		.PKT_TRANS_WRITE           (67),
		.PKT_TRANS_READ            (68),
		.PKT_TRANS_LOCK            (69),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (74),
		.PKT_BYTE_CNT_H            (73),
		.PKT_BYTE_CNT_L            (71),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                              //       clk_reset.reset
		.m0_address              (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src9_ready),                                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src9_valid),                                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src9_data),                                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src9_startofpacket),                                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src9_endofpacket),                                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src9_channel),                                                                             //                .channel
		.rf_sink_ready           (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                              // clk_reset.reset
		.in_data           (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                                        // (terminated)
		.csr_readdata      (),                                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                        // (terminated)
		.almost_full_data  (),                                                                                                            // (terminated)
		.almost_empty_data (),                                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                                        // (terminated)
		.out_empty         (),                                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                                        // (terminated)
		.out_error         (),                                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                                        // (terminated)
		.out_channel       ()                                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (64),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (65),
		.PKT_TRANS_POSTED          (66),
		.PKT_TRANS_WRITE           (67),
		.PKT_TRANS_READ            (68),
		.PKT_TRANS_LOCK            (69),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (74),
		.PKT_BYTE_CNT_H            (73),
		.PKT_BYTE_CNT_L            (71),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                //       clk_reset.reset
		.m0_address              (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src10_ready),                                                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src10_valid),                                                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src10_data),                                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src10_startofpacket),                                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src10_endofpacket),                                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src10_channel),                                                                              //                .channel
		.rf_sink_ready           (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                // clk_reset.reset
		.in_data           (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                                          // (terminated)
		.csr_readdata      (),                                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                          // (terminated)
		.almost_full_data  (),                                                                                                              // (terminated)
		.almost_empty_data (),                                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                                          // (terminated)
		.out_empty         (),                                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                                          // (terminated)
		.out_error         (),                                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                                          // (terminated)
		.out_channel       ()                                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (64),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (65),
		.PKT_TRANS_POSTED          (66),
		.PKT_TRANS_WRITE           (67),
		.PKT_TRANS_READ            (68),
		.PKT_TRANS_LOCK            (69),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (74),
		.PKT_BYTE_CNT_H            (73),
		.PKT_BYTE_CNT_L            (71),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                //       clk_reset.reset
		.m0_address              (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src11_ready),                                                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src11_valid),                                                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src11_data),                                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src11_startofpacket),                                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src11_endofpacket),                                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src11_channel),                                                                              //                .channel
		.rf_sink_ready           (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                // clk_reset.reset
		.in_data           (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                                          // (terminated)
		.csr_readdata      (),                                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                          // (terminated)
		.almost_full_data  (),                                                                                                              // (terminated)
		.almost_empty_data (),                                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                                          // (terminated)
		.out_empty         (),                                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                                          // (terminated)
		.out_error         (),                                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                                          // (terminated)
		.out_channel       ()                                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (64),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (65),
		.PKT_TRANS_POSTED          (66),
		.PKT_TRANS_WRITE           (67),
		.PKT_TRANS_READ            (68),
		.PKT_TRANS_LOCK            (69),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (74),
		.PKT_BYTE_CNT_H            (73),
		.PKT_BYTE_CNT_L            (71),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src12_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src12_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src12_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src12_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src12_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src12_channel),                                                                    //                .channel
		.rf_sink_ready           (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (64),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (65),
		.PKT_TRANS_POSTED          (66),
		.PKT_TRANS_WRITE           (67),
		.PKT_TRANS_READ            (68),
		.PKT_TRANS_LOCK            (69),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (74),
		.PKT_BYTE_CNT_H            (73),
		.PKT_BYTE_CNT_L            (71),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src13_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src13_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_001_src13_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src13_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src13_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src13_channel),                                                           //                .channel
		.rf_sink_ready           (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	nios_system_addr_router addr_router (
		.sink_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                              //       src.ready
		.src_valid          (addr_router_src_valid),                                                              //          .valid
		.src_data           (addr_router_src_data),                                                               //          .data
		.src_channel        (addr_router_src_channel),                                                            //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                         //          .endofpacket
	);

	nios_system_addr_router_001 addr_router_001 (
		.sink_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                   //          .valid
		.src_data           (addr_router_001_src_data),                                                    //          .data
		.src_channel        (addr_router_001_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                              //          .endofpacket
	);

	nios_system_id_router id_router (
		.sink_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                              //       src.ready
		.src_valid          (id_router_src_valid),                                                              //          .valid
		.src_data           (id_router_src_data),                                                               //          .data
		.src_channel        (id_router_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                         //          .endofpacket
	);

	nios_system_id_router_001 id_router_001 (
		.sink_ready         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                     //       src.ready
		.src_valid          (id_router_001_src_valid),                                                     //          .valid
		.src_data           (id_router_001_src_data),                                                      //          .data
		.src_channel        (id_router_001_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                //          .endofpacket
	);

	nios_system_id_router_002 id_router_002 (
		.sink_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                             //       src.ready
		.src_valid          (id_router_002_src_valid),                                             //          .valid
		.src_data           (id_router_002_src_data),                                              //          .data
		.src_channel        (id_router_002_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                        //          .endofpacket
	);

	nios_system_id_router_001 id_router_003 (
		.sink_ready         (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory_sram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                          //       src.ready
		.src_valid          (id_router_003_src_valid),                                                          //          .valid
		.src_data           (id_router_003_src_data),                                                           //          .data
		.src_channel        (id_router_003_src_channel),                                                        //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                     //          .endofpacket
	);

	nios_system_id_router_004 id_router_004 (
		.sink_ready         (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                     //       src.ready
		.src_valid          (id_router_004_src_valid),                                                     //          .valid
		.src_data           (id_router_004_src_data),                                                      //          .data
		.src_channel        (id_router_004_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                //          .endofpacket
	);

	nios_system_id_router_004 id_router_005 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                //          .valid
		.src_data           (id_router_005_src_data),                                                                 //          .data
		.src_channel        (id_router_005_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                           //          .endofpacket
	);

	nios_system_id_router_004 id_router_006 (
		.sink_ready         (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                      //       src.ready
		.src_valid          (id_router_006_src_valid),                                                      //          .valid
		.src_data           (id_router_006_src_data),                                                       //          .data
		.src_channel        (id_router_006_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                 //          .endofpacket
	);

	nios_system_id_router_004 id_router_007 (
		.sink_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                        //       src.ready
		.src_valid          (id_router_007_src_valid),                                                        //          .valid
		.src_data           (id_router_007_src_data),                                                         //          .data
		.src_channel        (id_router_007_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                   //          .endofpacket
	);

	nios_system_id_router_004 id_router_008 (
		.sink_ready         (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                                          //       src.ready
		.src_valid          (id_router_008_src_valid),                                                                          //          .valid
		.src_data           (id_router_008_src_data),                                                                           //          .data
		.src_channel        (id_router_008_src_channel),                                                                        //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                                  //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                                     //          .endofpacket
	);

	nios_system_id_router_004 id_router_009 (
		.sink_ready         (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                                         //       src.ready
		.src_valid          (id_router_009_src_valid),                                                                         //          .valid
		.src_data           (id_router_009_src_data),                                                                          //          .data
		.src_channel        (id_router_009_src_channel),                                                                       //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                                 //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                                    //          .endofpacket
	);

	nios_system_id_router_004 id_router_010 (
		.sink_ready         (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                        // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                                               //       src.ready
		.src_valid          (id_router_010_src_valid),                                                                               //          .valid
		.src_data           (id_router_010_src_data),                                                                                //          .data
		.src_channel        (id_router_010_src_channel),                                                                             //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                                                       //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                                          //          .endofpacket
	);

	nios_system_id_router_004 id_router_011 (
		.sink_ready         (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                    // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                                           //       src.ready
		.src_valid          (id_router_011_src_valid),                                                                           //          .valid
		.src_data           (id_router_011_src_data),                                                                            //          .data
		.src_channel        (id_router_011_src_channel),                                                                         //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                                                   //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                                      //          .endofpacket
	);

	nios_system_id_router_004 id_router_012 (
		.sink_ready         (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (expansion_jp1_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                                             //       src.ready
		.src_valid          (id_router_012_src_valid),                                                                             //          .valid
		.src_data           (id_router_012_src_data),                                                                              //          .data
		.src_channel        (id_router_012_src_channel),                                                                           //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                                                     //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                                                        //          .endofpacket
	);

	nios_system_id_router_004 id_router_013 (
		.sink_ready         (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (expansion_jp2_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                                             //       src.ready
		.src_valid          (id_router_013_src_valid),                                                                             //          .valid
		.src_data           (id_router_013_src_data),                                                                              //          .data
		.src_channel        (id_router_013_src_channel),                                                                           //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                                                     //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                                                        //          .endofpacket
	);

	nios_system_id_router_004 id_router_014 (
		.sink_ready         (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_014_src_valid),                                                                   //          .valid
		.src_data           (id_router_014_src_data),                                                                    //          .data
		.src_channel        (id_router_014_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                                              //          .endofpacket
	);

	nios_system_id_router_004 id_router_015 (
		.sink_ready         (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory_sram_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                                          //       src.ready
		.src_valid          (id_router_015_src_valid),                                                          //          .valid
		.src_data           (id_router_015_src_data),                                                           //          .data
		.src_channel        (id_router_015_src_channel),                                                        //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                                     //          .endofpacket
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (46),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (66),
		.PKT_BYTE_CNT_H            (55),
		.PKT_BYTE_CNT_L            (53),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (61),
		.PKT_BURST_SIZE_L          (59),
		.PKT_BURST_TYPE_H          (63),
		.PKT_BURST_TYPE_L          (62),
		.PKT_BURSTWRAP_H           (58),
		.PKT_BURSTWRAP_L           (56),
		.PKT_TRANS_COMPRESSED_READ (47),
		.PKT_TRANS_WRITE           (49),
		.PKT_TRANS_READ            (50),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (86),
		.ST_CHANNEL_W              (16),
		.OUT_BYTE_CNT_H            (54),
		.OUT_BURSTWRAP_H           (58),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_n),                          // reset_in0.reset
		.reset_in1  (cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk),                               //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_in2  (1'b0),                              // (terminated)
		.reset_in3  (1'b0),                              // (terminated)
		.reset_in4  (1'b0),                              // (terminated)
		.reset_in5  (1'b0),                              // (terminated)
		.reset_in6  (1'b0),                              // (terminated)
		.reset_in7  (1'b0),                              // (terminated)
		.reset_in8  (1'b0),                              // (terminated)
		.reset_in9  (1'b0),                              // (terminated)
		.reset_in10 (1'b0),                              // (terminated)
		.reset_in11 (1'b0),                              // (terminated)
		.reset_in12 (1'b0),                              // (terminated)
		.reset_in13 (1'b0),                              // (terminated)
		.reset_in14 (1'b0),                              // (terminated)
		.reset_in15 (1'b0)                               // (terminated)
	);

	nios_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (clk),                                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_001_src_ready),              //      sink.ready
		.sink_channel        (addr_router_001_src_channel),            //          .channel
		.sink_data           (addr_router_001_src_data),               //          .data
		.sink_startofpacket  (addr_router_001_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_001_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_001_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk),                                   //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (clk),                                   //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_001 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_003 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_004 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_005 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_006 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_007 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_008 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_009 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_010 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_011 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_012 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_013 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_014 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_015 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk),                                   //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (clk),                                   //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_002_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_004_src0_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_005_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_006_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_007_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_008_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_009_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_010_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_010_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_011_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_011_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_012_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_013_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_014_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_015_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (64),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (73),
		.IN_PKT_BYTE_CNT_L             (71),
		.IN_PKT_TRANS_COMPRESSED_READ  (65),
		.IN_PKT_BURSTWRAP_H            (76),
		.IN_PKT_BURSTWRAP_L            (74),
		.IN_PKT_BURST_SIZE_H           (79),
		.IN_PKT_BURST_SIZE_L           (77),
		.IN_PKT_RESPONSE_STATUS_H      (103),
		.IN_PKT_RESPONSE_STATUS_L      (102),
		.IN_PKT_TRANS_EXCLUSIVE        (70),
		.IN_PKT_BURST_TYPE_H           (81),
		.IN_PKT_BURST_TYPE_L           (80),
		.IN_ST_DATA_W                  (104),
		.OUT_PKT_ADDR_H                (46),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (55),
		.OUT_PKT_BYTE_CNT_L            (53),
		.OUT_PKT_TRANS_COMPRESSED_READ (47),
		.OUT_PKT_BURST_SIZE_H          (61),
		.OUT_PKT_BURST_SIZE_L          (59),
		.OUT_PKT_RESPONSE_STATUS_H     (85),
		.OUT_PKT_RESPONSE_STATUS_L     (84),
		.OUT_PKT_TRANS_EXCLUSIVE       (52),
		.OUT_PKT_BURST_TYPE_H          (63),
		.OUT_PKT_BURST_TYPE_L          (62),
		.OUT_ST_DATA_W                 (86),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (clk),                                //       clk.clk
		.reset                (rst_controller_reset_out_reset),     // clk_reset.reset
		.in_valid             (cmd_xbar_mux_002_src_valid),         //      sink.valid
		.in_channel           (cmd_xbar_mux_002_src_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_mux_002_src_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_002_src_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_mux_002_src_ready),         //          .ready
		.in_data              (cmd_xbar_mux_002_src_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (46),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (55),
		.IN_PKT_BYTE_CNT_L             (53),
		.IN_PKT_TRANS_COMPRESSED_READ  (47),
		.IN_PKT_BURSTWRAP_H            (58),
		.IN_PKT_BURSTWRAP_L            (56),
		.IN_PKT_BURST_SIZE_H           (61),
		.IN_PKT_BURST_SIZE_L           (59),
		.IN_PKT_RESPONSE_STATUS_H      (85),
		.IN_PKT_RESPONSE_STATUS_L      (84),
		.IN_PKT_TRANS_EXCLUSIVE        (52),
		.IN_PKT_BURST_TYPE_H           (63),
		.IN_PKT_BURST_TYPE_L           (62),
		.IN_ST_DATA_W                  (86),
		.OUT_PKT_ADDR_H                (64),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (73),
		.OUT_PKT_BYTE_CNT_L            (71),
		.OUT_PKT_TRANS_COMPRESSED_READ (65),
		.OUT_PKT_BURST_SIZE_H          (79),
		.OUT_PKT_BURST_SIZE_L          (77),
		.OUT_PKT_RESPONSE_STATUS_H     (103),
		.OUT_PKT_RESPONSE_STATUS_L     (102),
		.OUT_PKT_TRANS_EXCLUSIVE       (70),
		.OUT_PKT_BURST_TYPE_H          (81),
		.OUT_PKT_BURST_TYPE_L          (80),
		.OUT_ST_DATA_W                 (104),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_001 (
		.clk                  (clk),                                 //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_002_src_valid),             //      sink.valid
		.in_channel           (id_router_002_src_channel),           //          .channel
		.in_startofpacket     (id_router_002_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_002_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_002_src_ready),             //          .ready
		.in_data              (id_router_002_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clk),                            //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

endmodule

// nios_system.v

// Generated using ACDS version 13.1 162 at 2018.04.13.21:38:49

`timescale 1 ps / 1 ps
module nios_system (
		input  wire        reset_n,                              //                   clk_clk_in_reset.reset_n
		inout  wire [31:0] GPIO_0_to_and_from_the_Expansion_JP1, //   Expansion_JP1_external_interface.export
		output wire [9:0]  LEDG_from_the_Green_LEDs,             //      Green_LEDs_external_interface.export
		output wire [11:0] zs_addr_from_the_sdram,               //                         sdram_wire.addr
		output wire [1:0]  zs_ba_from_the_sdram,                 //                                   .ba
		output wire        zs_cas_n_from_the_sdram,              //                                   .cas_n
		output wire        zs_cke_from_the_sdram,                //                                   .cke
		output wire        zs_cs_n_from_the_sdram,               //                                   .cs_n
		inout  wire [15:0] zs_dq_to_and_from_the_sdram,          //                                   .dq
		output wire [1:0]  zs_dqm_from_the_sdram,                //                                   .dqm
		output wire        zs_ras_n_from_the_sdram,              //                                   .ras_n
		output wire        zs_we_n_from_the_sdram,               //                                   .we_n
		inout  wire [31:0] GPIO_1_to_and_from_the_Expansion_JP2, //   Expansion_JP2_external_interface.export
		input  wire        UART_RXD_to_the_Serial_port,          //     Serial_port_external_interface.RXD
		output wire        UART_TXD_from_the_Serial_port,        //                                   .TXD
		input  wire        clk,                                  //                         clk_clk_in.clk
		input  wire [2:0]  KEY_to_the_Pushbuttons,               //     Pushbuttons_external_interface.export
		input  wire [9:0]  SW_to_the_Slider_switches,            // Slider_switches_external_interface.export
		output wire [7:0]  HEX0_from_the_HEX3_HEX0,              //       HEX3_HEX0_external_interface.HEX0
		output wire [7:0]  HEX1_from_the_HEX3_HEX0,              //                                   .HEX1
		output wire [7:0]  HEX2_from_the_HEX3_HEX0,              //                                   .HEX2
		output wire [7:0]  HEX3_from_the_HEX3_HEX0               //                                   .HEX3
	);

	wire  [15:0] mm_interconnect_0_interval_timer_s1_writedata;                           // mm_interconnect_0:Interval_timer_s1_writedata -> Interval_timer:writedata
	wire   [2:0] mm_interconnect_0_interval_timer_s1_address;                             // mm_interconnect_0:Interval_timer_s1_address -> Interval_timer:address
	wire         mm_interconnect_0_interval_timer_s1_chipselect;                          // mm_interconnect_0:Interval_timer_s1_chipselect -> Interval_timer:chipselect
	wire         mm_interconnect_0_interval_timer_s1_write;                               // mm_interconnect_0:Interval_timer_s1_write -> Interval_timer:write_n
	wire  [15:0] mm_interconnect_0_interval_timer_s1_readdata;                            // Interval_timer:readdata -> mm_interconnect_0:Interval_timer_s1_readdata
	wire  [31:0] mm_interconnect_0_slider_switches_avalon_parallel_port_slave_writedata;  // mm_interconnect_0:Slider_switches_avalon_parallel_port_slave_writedata -> Slider_switches:writedata
	wire   [1:0] mm_interconnect_0_slider_switches_avalon_parallel_port_slave_address;    // mm_interconnect_0:Slider_switches_avalon_parallel_port_slave_address -> Slider_switches:address
	wire         mm_interconnect_0_slider_switches_avalon_parallel_port_slave_chipselect; // mm_interconnect_0:Slider_switches_avalon_parallel_port_slave_chipselect -> Slider_switches:chipselect
	wire         mm_interconnect_0_slider_switches_avalon_parallel_port_slave_write;      // mm_interconnect_0:Slider_switches_avalon_parallel_port_slave_write -> Slider_switches:write
	wire         mm_interconnect_0_slider_switches_avalon_parallel_port_slave_read;       // mm_interconnect_0:Slider_switches_avalon_parallel_port_slave_read -> Slider_switches:read
	wire  [31:0] mm_interconnect_0_slider_switches_avalon_parallel_port_slave_readdata;   // Slider_switches:readdata -> mm_interconnect_0:Slider_switches_avalon_parallel_port_slave_readdata
	wire   [3:0] mm_interconnect_0_slider_switches_avalon_parallel_port_slave_byteenable; // mm_interconnect_0:Slider_switches_avalon_parallel_port_slave_byteenable -> Slider_switches:byteenable
	wire  [31:0] mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_writedata;      // mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_writedata -> Pushbuttons:writedata
	wire   [1:0] mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_address;        // mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_address -> Pushbuttons:address
	wire         mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_chipselect;     // mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_chipselect -> Pushbuttons:chipselect
	wire         mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_write;          // mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_write -> Pushbuttons:write
	wire         mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_read;           // mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_read -> Pushbuttons:read
	wire  [31:0] mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_readdata;       // Pushbuttons:readdata -> mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_readdata
	wire   [3:0] mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_byteenable;     // mm_interconnect_0:Pushbuttons_avalon_parallel_port_slave_byteenable -> Pushbuttons:byteenable
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                           // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                          // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire         cpu_data_master_waitrequest;                                             // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                               // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [28:0] cpu_data_master_address;                                                 // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire         cpu_data_master_write;                                                   // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire         cpu_data_master_read;                                                    // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                                // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_debugaccess;                                             // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire   [3:0] cpu_data_master_byteenable;                                              // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                            // mm_interconnect_0:Onchip_memory_s1_writedata -> Onchip_memory:writedata
	wire  [10:0] mm_interconnect_0_onchip_memory_s1_address;                              // mm_interconnect_0:Onchip_memory_s1_address -> Onchip_memory:address
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                           // mm_interconnect_0:Onchip_memory_s1_chipselect -> Onchip_memory:chipselect
	wire         mm_interconnect_0_onchip_memory_s1_clken;                                // mm_interconnect_0:Onchip_memory_s1_clken -> Onchip_memory:clken
	wire         mm_interconnect_0_onchip_memory_s1_write;                                // mm_interconnect_0:Onchip_memory_s1_write -> Onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                             // Onchip_memory:readdata -> mm_interconnect_0:Onchip_memory_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                           // mm_interconnect_0:Onchip_memory_s1_byteenable -> Onchip_memory:byteenable
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                  // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                    // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [21:0] mm_interconnect_0_sdram_s1_address;                                      // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                                   // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                                        // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                                         // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                     // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                   // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;                     // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;                       // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;                         // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;                           // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                            // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;                        // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;                     // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;                      // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire         cpu_instruction_master_waitrequest;                                      // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                                          // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                             // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                                         // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;               // JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                 // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                   // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                     // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> JTAG_UART:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                      // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> JTAG_UART:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                  // JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_serial_port_avalon_rs232_slave_writedata;              // mm_interconnect_0:Serial_port_avalon_rs232_slave_writedata -> Serial_port:writedata
	wire   [0:0] mm_interconnect_0_serial_port_avalon_rs232_slave_address;                // mm_interconnect_0:Serial_port_avalon_rs232_slave_address -> Serial_port:address
	wire         mm_interconnect_0_serial_port_avalon_rs232_slave_chipselect;             // mm_interconnect_0:Serial_port_avalon_rs232_slave_chipselect -> Serial_port:chipselect
	wire         mm_interconnect_0_serial_port_avalon_rs232_slave_write;                  // mm_interconnect_0:Serial_port_avalon_rs232_slave_write -> Serial_port:write
	wire         mm_interconnect_0_serial_port_avalon_rs232_slave_read;                   // mm_interconnect_0:Serial_port_avalon_rs232_slave_read -> Serial_port:read
	wire  [31:0] mm_interconnect_0_serial_port_avalon_rs232_slave_readdata;               // Serial_port:readdata -> mm_interconnect_0:Serial_port_avalon_rs232_slave_readdata
	wire   [3:0] mm_interconnect_0_serial_port_avalon_rs232_slave_byteenable;             // mm_interconnect_0:Serial_port_avalon_rs232_slave_byteenable -> Serial_port:byteenable
	wire  [31:0] mm_interconnect_0_onchip_memory_s2_writedata;                            // mm_interconnect_0:Onchip_memory_s2_writedata -> Onchip_memory:writedata2
	wire  [10:0] mm_interconnect_0_onchip_memory_s2_address;                              // mm_interconnect_0:Onchip_memory_s2_address -> Onchip_memory:address2
	wire         mm_interconnect_0_onchip_memory_s2_chipselect;                           // mm_interconnect_0:Onchip_memory_s2_chipselect -> Onchip_memory:chipselect2
	wire         mm_interconnect_0_onchip_memory_s2_clken;                                // mm_interconnect_0:Onchip_memory_s2_clken -> Onchip_memory:clken2
	wire         mm_interconnect_0_onchip_memory_s2_write;                                // mm_interconnect_0:Onchip_memory_s2_write -> Onchip_memory:write2
	wire  [31:0] mm_interconnect_0_onchip_memory_s2_readdata;                             // Onchip_memory:readdata2 -> mm_interconnect_0:Onchip_memory_s2_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory_s2_byteenable;                           // mm_interconnect_0:Onchip_memory_s2_byteenable -> Onchip_memory:byteenable2
	wire  [31:0] mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_writedata;    // mm_interconnect_0:Expansion_JP1_avalon_parallel_port_slave_writedata -> Expansion_JP1:writedata
	wire   [1:0] mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_address;      // mm_interconnect_0:Expansion_JP1_avalon_parallel_port_slave_address -> Expansion_JP1:address
	wire         mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_chipselect;   // mm_interconnect_0:Expansion_JP1_avalon_parallel_port_slave_chipselect -> Expansion_JP1:chipselect
	wire         mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_write;        // mm_interconnect_0:Expansion_JP1_avalon_parallel_port_slave_write -> Expansion_JP1:write
	wire         mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_read;         // mm_interconnect_0:Expansion_JP1_avalon_parallel_port_slave_read -> Expansion_JP1:read
	wire  [31:0] mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_readdata;     // Expansion_JP1:readdata -> mm_interconnect_0:Expansion_JP1_avalon_parallel_port_slave_readdata
	wire   [3:0] mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_byteenable;   // mm_interconnect_0:Expansion_JP1_avalon_parallel_port_slave_byteenable -> Expansion_JP1:byteenable
	wire  [31:0] mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_writedata;    // mm_interconnect_0:Expansion_JP2_avalon_parallel_port_slave_writedata -> Expansion_JP2:writedata
	wire   [1:0] mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_address;      // mm_interconnect_0:Expansion_JP2_avalon_parallel_port_slave_address -> Expansion_JP2:address
	wire         mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_chipselect;   // mm_interconnect_0:Expansion_JP2_avalon_parallel_port_slave_chipselect -> Expansion_JP2:chipselect
	wire         mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_write;        // mm_interconnect_0:Expansion_JP2_avalon_parallel_port_slave_write -> Expansion_JP2:write
	wire         mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_read;         // mm_interconnect_0:Expansion_JP2_avalon_parallel_port_slave_read -> Expansion_JP2:read
	wire  [31:0] mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_readdata;     // Expansion_JP2:readdata -> mm_interconnect_0:Expansion_JP2_avalon_parallel_port_slave_readdata
	wire   [3:0] mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_byteenable;   // mm_interconnect_0:Expansion_JP2_avalon_parallel_port_slave_byteenable -> Expansion_JP2:byteenable
	wire  [31:0] mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_writedata;        // mm_interconnect_0:HEX3_HEX0_avalon_parallel_port_slave_writedata -> HEX3_HEX0:writedata
	wire   [1:0] mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_address;          // mm_interconnect_0:HEX3_HEX0_avalon_parallel_port_slave_address -> HEX3_HEX0:address
	wire         mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_chipselect;       // mm_interconnect_0:HEX3_HEX0_avalon_parallel_port_slave_chipselect -> HEX3_HEX0:chipselect
	wire         mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_write;            // mm_interconnect_0:HEX3_HEX0_avalon_parallel_port_slave_write -> HEX3_HEX0:write
	wire         mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_read;             // mm_interconnect_0:HEX3_HEX0_avalon_parallel_port_slave_read -> HEX3_HEX0:read
	wire  [31:0] mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_readdata;         // HEX3_HEX0:readdata -> mm_interconnect_0:HEX3_HEX0_avalon_parallel_port_slave_readdata
	wire   [3:0] mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_byteenable;       // mm_interconnect_0:HEX3_HEX0_avalon_parallel_port_slave_byteenable -> HEX3_HEX0:byteenable
	wire  [31:0] mm_interconnect_0_onchip_memory_sram_s2_writedata;                       // mm_interconnect_0:Onchip_memory_SRAM_s2_writedata -> Onchip_memory_SRAM:writedata2
	wire  [10:0] mm_interconnect_0_onchip_memory_sram_s2_address;                         // mm_interconnect_0:Onchip_memory_SRAM_s2_address -> Onchip_memory_SRAM:address2
	wire         mm_interconnect_0_onchip_memory_sram_s2_chipselect;                      // mm_interconnect_0:Onchip_memory_SRAM_s2_chipselect -> Onchip_memory_SRAM:chipselect2
	wire         mm_interconnect_0_onchip_memory_sram_s2_clken;                           // mm_interconnect_0:Onchip_memory_SRAM_s2_clken -> Onchip_memory_SRAM:clken2
	wire         mm_interconnect_0_onchip_memory_sram_s2_write;                           // mm_interconnect_0:Onchip_memory_SRAM_s2_write -> Onchip_memory_SRAM:write2
	wire  [31:0] mm_interconnect_0_onchip_memory_sram_s2_readdata;                        // Onchip_memory_SRAM:readdata2 -> mm_interconnect_0:Onchip_memory_SRAM_s2_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory_sram_s2_byteenable;                      // mm_interconnect_0:Onchip_memory_SRAM_s2_byteenable -> Onchip_memory_SRAM:byteenable2
	wire  [31:0] mm_interconnect_0_onchip_memory_sram_s1_writedata;                       // mm_interconnect_0:Onchip_memory_SRAM_s1_writedata -> Onchip_memory_SRAM:writedata
	wire  [10:0] mm_interconnect_0_onchip_memory_sram_s1_address;                         // mm_interconnect_0:Onchip_memory_SRAM_s1_address -> Onchip_memory_SRAM:address
	wire         mm_interconnect_0_onchip_memory_sram_s1_chipselect;                      // mm_interconnect_0:Onchip_memory_SRAM_s1_chipselect -> Onchip_memory_SRAM:chipselect
	wire         mm_interconnect_0_onchip_memory_sram_s1_clken;                           // mm_interconnect_0:Onchip_memory_SRAM_s1_clken -> Onchip_memory_SRAM:clken
	wire         mm_interconnect_0_onchip_memory_sram_s1_write;                           // mm_interconnect_0:Onchip_memory_SRAM_s1_write -> Onchip_memory_SRAM:write
	wire  [31:0] mm_interconnect_0_onchip_memory_sram_s1_readdata;                        // Onchip_memory_SRAM:readdata -> mm_interconnect_0:Onchip_memory_SRAM_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory_sram_s1_byteenable;                      // mm_interconnect_0:Onchip_memory_SRAM_s1_byteenable -> Onchip_memory_SRAM:byteenable
	wire  [31:0] mm_interconnect_0_green_leds_avalon_parallel_port_slave_writedata;       // mm_interconnect_0:Green_LEDs_avalon_parallel_port_slave_writedata -> Green_LEDs:writedata
	wire   [1:0] mm_interconnect_0_green_leds_avalon_parallel_port_slave_address;         // mm_interconnect_0:Green_LEDs_avalon_parallel_port_slave_address -> Green_LEDs:address
	wire         mm_interconnect_0_green_leds_avalon_parallel_port_slave_chipselect;      // mm_interconnect_0:Green_LEDs_avalon_parallel_port_slave_chipselect -> Green_LEDs:chipselect
	wire         mm_interconnect_0_green_leds_avalon_parallel_port_slave_write;           // mm_interconnect_0:Green_LEDs_avalon_parallel_port_slave_write -> Green_LEDs:write
	wire         mm_interconnect_0_green_leds_avalon_parallel_port_slave_read;            // mm_interconnect_0:Green_LEDs_avalon_parallel_port_slave_read -> Green_LEDs:read
	wire  [31:0] mm_interconnect_0_green_leds_avalon_parallel_port_slave_readdata;        // Green_LEDs:readdata -> mm_interconnect_0:Green_LEDs_avalon_parallel_port_slave_readdata
	wire   [3:0] mm_interconnect_0_green_leds_avalon_parallel_port_slave_byteenable;      // mm_interconnect_0:Green_LEDs_avalon_parallel_port_slave_byteenable -> Green_LEDs:byteenable
	wire         irq_mapper_receiver0_irq;                                                // JTAG_UART:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                // Interval_timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                // Serial_port:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                // Pushbuttons:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                // Expansion_JP1:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                                // Expansion_JP2:irq -> irq_mapper:receiver5_irq
	wire  [31:0] cpu_d_irq_irq;                                                           // irq_mapper:sender_irq -> cpu:d_irq
	wire         rst_controller_reset_out_reset;                                          // rst_controller:reset_out -> [Expansion_JP1:reset, Expansion_JP2:reset, Green_LEDs:reset, HEX3_HEX0:reset, Interval_timer:reset_n, JTAG_UART:rst_n, Onchip_memory:reset, Onchip_memory:reset2, Onchip_memory_SRAM:reset, Onchip_memory_SRAM:reset2, Pushbuttons:reset, Serial_port:reset, Slider_switches:reset, cpu:reset_n, irq_mapper:reset, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram:reset_n, sysid:reset_n]
	wire         rst_controller_reset_out_reset_req;                                      // rst_controller:reset_req -> [Onchip_memory:reset_req, Onchip_memory:reset_req2, Onchip_memory_SRAM:reset_req, Onchip_memory_SRAM:reset_req2, cpu:reset_req, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                                       // cpu:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	nios_system_Onchip_memory onchip_memory (
		.clk         (clk),                                           //   clk1.clk
		.address     (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata    (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),            //       .reset_req
		.address2    (mm_interconnect_0_onchip_memory_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_onchip_memory_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_onchip_memory_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_onchip_memory_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_onchip_memory_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_onchip_memory_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_onchip_memory_s2_byteenable), //       .byteenable
		.clk2        (clk),                                           //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),                // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req)             //       .reset_req
	);

	nios_system_JTAG_UART jtag_uart (
		.clk            (clk),                                                       //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	nios_system_Interval_timer interval_timer (
		.clk        (clk),                                            //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                // reset.reset_n
		.address    (mm_interconnect_0_interval_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_interval_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_interval_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_interval_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_interval_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                        //   irq.irq
	);

	nios_system_sdram sdram (
		.clk            (clk),                                      //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (zs_addr_from_the_sdram),                   //  wire.export
		.zs_ba          (zs_ba_from_the_sdram),                     //      .export
		.zs_cas_n       (zs_cas_n_from_the_sdram),                  //      .export
		.zs_cke         (zs_cke_from_the_sdram),                    //      .export
		.zs_cs_n        (zs_cs_n_from_the_sdram),                   //      .export
		.zs_dq          (zs_dq_to_and_from_the_sdram),              //      .export
		.zs_dqm         (zs_dqm_from_the_sdram),                    //      .export
		.zs_ras_n       (zs_ras_n_from_the_sdram),                  //      .export
		.zs_we_n        (zs_we_n_from_the_sdram)                    //      .export
	);

	nios_system_Green_LEDs green_leds (
		.clk        (clk),                                                                //                clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                     //          clock_reset_reset.reset
		.address    (mm_interconnect_0_green_leds_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_green_leds_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_green_leds_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_green_leds_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_green_leds_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_green_leds_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_green_leds_avalon_parallel_port_slave_readdata),   //                           .readdata
		.LEDG       (LEDG_from_the_Green_LEDs)                                            //         external_interface.export
	);

	nios_system_HEX3_HEX0 hex3_hex0 (
		.clk        (clk),                                                               //                clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                    //          clock_reset_reset.reset
		.address    (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_readdata),   //                           .readdata
		.HEX0       (HEX0_from_the_HEX3_HEX0),                                           //         external_interface.export
		.HEX1       (HEX1_from_the_HEX3_HEX0),                                           //                           .export
		.HEX2       (HEX2_from_the_HEX3_HEX0),                                           //                           .export
		.HEX3       (HEX3_from_the_HEX3_HEX0)                                            //                           .export
	);

	nios_system_Slider_switches slider_switches (
		.clk        (clk),                                                                     //                clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                          //          clock_reset_reset.reset
		.address    (mm_interconnect_0_slider_switches_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_slider_switches_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_slider_switches_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_slider_switches_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_slider_switches_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_slider_switches_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_slider_switches_avalon_parallel_port_slave_readdata),   //                           .readdata
		.SW         (SW_to_the_Slider_switches)                                                //         external_interface.export
	);

	nios_system_Pushbuttons pushbuttons (
		.clk        (clk),                                                                 //                clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                      //          clock_reset_reset.reset
		.address    (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_readdata),   //                           .readdata
		.KEY        (KEY_to_the_Pushbuttons),                                              //         external_interface.export
		.irq        (irq_mapper_receiver3_irq)                                             //                  interrupt.irq
	);

	nios_system_Expansion_JP1 expansion_jp1 (
		.clk        (clk),                                                                   //                clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                        //          clock_reset_reset.reset
		.address    (mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_readdata),   //                           .readdata
		.GPIO_0     (GPIO_0_to_and_from_the_Expansion_JP1),                                  //         external_interface.export
		.irq        (irq_mapper_receiver4_irq)                                               //                  interrupt.irq
	);

	nios_system_Expansion_JP2 expansion_jp2 (
		.clk        (clk),                                                                   //                clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                        //          clock_reset_reset.reset
		.address    (mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_readdata),   //                           .readdata
		.GPIO_1     (GPIO_1_to_and_from_the_Expansion_JP2),                                  //         external_interface.export
		.irq        (irq_mapper_receiver5_irq)                                               //                  interrupt.irq
	);

	nios_system_Serial_port serial_port (
		.clk        (clk),                                                         //        clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                              //  clock_reset_reset.reset
		.address    (mm_interconnect_0_serial_port_avalon_rs232_slave_address),    // avalon_rs232_slave.address
		.chipselect (mm_interconnect_0_serial_port_avalon_rs232_slave_chipselect), //                   .chipselect
		.byteenable (mm_interconnect_0_serial_port_avalon_rs232_slave_byteenable), //                   .byteenable
		.read       (mm_interconnect_0_serial_port_avalon_rs232_slave_read),       //                   .read
		.write      (mm_interconnect_0_serial_port_avalon_rs232_slave_write),      //                   .write
		.writedata  (mm_interconnect_0_serial_port_avalon_rs232_slave_writedata),  //                   .writedata
		.readdata   (mm_interconnect_0_serial_port_avalon_rs232_slave_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver2_irq),                                    //          interrupt.irq
		.UART_RXD   (UART_RXD_to_the_Serial_port),                                 // external_interface.export
		.UART_TXD   (UART_TXD_from_the_Serial_port)                                //                   .export
	);

	nios_system_Onchip_memory_SRAM onchip_memory_sram (
		.clk         (clk),                                                //   clk1.clk
		.address     (mm_interconnect_0_onchip_memory_sram_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_onchip_memory_sram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_onchip_memory_sram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_onchip_memory_sram_s1_write),      //       .write
		.readdata    (mm_interconnect_0_onchip_memory_sram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_onchip_memory_sram_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_onchip_memory_sram_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                     // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),                 //       .reset_req
		.address2    (mm_interconnect_0_onchip_memory_sram_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_onchip_memory_sram_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_onchip_memory_sram_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_onchip_memory_sram_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_onchip_memory_sram_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_onchip_memory_sram_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_onchip_memory_sram_s2_byteenable), //       .byteenable
		.clk2        (clk),                                                //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),                     // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req)                  //       .reset_req
	);

	nios_system_cpu cpu (
		.clk                                   (clk),                                                 //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	nios_system_sysid sysid (
		.clock    (clk),                                            //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                           (clk),                                                                     //                                    clk_clk.clk
		.cpu_reset_n_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                                          //          cpu_reset_n_reset_bridge_in_reset.reset
		.cpu_data_master_address                               (cpu_data_master_address),                                                 //                            cpu_data_master.address
		.cpu_data_master_waitrequest                           (cpu_data_master_waitrequest),                                             //                                           .waitrequest
		.cpu_data_master_byteenable                            (cpu_data_master_byteenable),                                              //                                           .byteenable
		.cpu_data_master_read                                  (cpu_data_master_read),                                                    //                                           .read
		.cpu_data_master_readdata                              (cpu_data_master_readdata),                                                //                                           .readdata
		.cpu_data_master_write                                 (cpu_data_master_write),                                                   //                                           .write
		.cpu_data_master_writedata                             (cpu_data_master_writedata),                                               //                                           .writedata
		.cpu_data_master_debugaccess                           (cpu_data_master_debugaccess),                                             //                                           .debugaccess
		.cpu_instruction_master_address                        (cpu_instruction_master_address),                                          //                     cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                    (cpu_instruction_master_waitrequest),                                      //                                           .waitrequest
		.cpu_instruction_master_read                           (cpu_instruction_master_read),                                             //                                           .read
		.cpu_instruction_master_readdata                       (cpu_instruction_master_readdata),                                         //                                           .readdata
		.cpu_jtag_debug_module_address                         (mm_interconnect_0_cpu_jtag_debug_module_address),                         //                      cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write                           (mm_interconnect_0_cpu_jtag_debug_module_write),                           //                                           .write
		.cpu_jtag_debug_module_read                            (mm_interconnect_0_cpu_jtag_debug_module_read),                            //                                           .read
		.cpu_jtag_debug_module_readdata                        (mm_interconnect_0_cpu_jtag_debug_module_readdata),                        //                                           .readdata
		.cpu_jtag_debug_module_writedata                       (mm_interconnect_0_cpu_jtag_debug_module_writedata),                       //                                           .writedata
		.cpu_jtag_debug_module_byteenable                      (mm_interconnect_0_cpu_jtag_debug_module_byteenable),                      //                                           .byteenable
		.cpu_jtag_debug_module_waitrequest                     (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),                     //                                           .waitrequest
		.cpu_jtag_debug_module_debugaccess                     (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),                     //                                           .debugaccess
		.Expansion_JP1_avalon_parallel_port_slave_address      (mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_address),      //   Expansion_JP1_avalon_parallel_port_slave.address
		.Expansion_JP1_avalon_parallel_port_slave_write        (mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_write),        //                                           .write
		.Expansion_JP1_avalon_parallel_port_slave_read         (mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_read),         //                                           .read
		.Expansion_JP1_avalon_parallel_port_slave_readdata     (mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_readdata),     //                                           .readdata
		.Expansion_JP1_avalon_parallel_port_slave_writedata    (mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_writedata),    //                                           .writedata
		.Expansion_JP1_avalon_parallel_port_slave_byteenable   (mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_byteenable),   //                                           .byteenable
		.Expansion_JP1_avalon_parallel_port_slave_chipselect   (mm_interconnect_0_expansion_jp1_avalon_parallel_port_slave_chipselect),   //                                           .chipselect
		.Expansion_JP2_avalon_parallel_port_slave_address      (mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_address),      //   Expansion_JP2_avalon_parallel_port_slave.address
		.Expansion_JP2_avalon_parallel_port_slave_write        (mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_write),        //                                           .write
		.Expansion_JP2_avalon_parallel_port_slave_read         (mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_read),         //                                           .read
		.Expansion_JP2_avalon_parallel_port_slave_readdata     (mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_readdata),     //                                           .readdata
		.Expansion_JP2_avalon_parallel_port_slave_writedata    (mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_writedata),    //                                           .writedata
		.Expansion_JP2_avalon_parallel_port_slave_byteenable   (mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_byteenable),   //                                           .byteenable
		.Expansion_JP2_avalon_parallel_port_slave_chipselect   (mm_interconnect_0_expansion_jp2_avalon_parallel_port_slave_chipselect),   //                                           .chipselect
		.Green_LEDs_avalon_parallel_port_slave_address         (mm_interconnect_0_green_leds_avalon_parallel_port_slave_address),         //      Green_LEDs_avalon_parallel_port_slave.address
		.Green_LEDs_avalon_parallel_port_slave_write           (mm_interconnect_0_green_leds_avalon_parallel_port_slave_write),           //                                           .write
		.Green_LEDs_avalon_parallel_port_slave_read            (mm_interconnect_0_green_leds_avalon_parallel_port_slave_read),            //                                           .read
		.Green_LEDs_avalon_parallel_port_slave_readdata        (mm_interconnect_0_green_leds_avalon_parallel_port_slave_readdata),        //                                           .readdata
		.Green_LEDs_avalon_parallel_port_slave_writedata       (mm_interconnect_0_green_leds_avalon_parallel_port_slave_writedata),       //                                           .writedata
		.Green_LEDs_avalon_parallel_port_slave_byteenable      (mm_interconnect_0_green_leds_avalon_parallel_port_slave_byteenable),      //                                           .byteenable
		.Green_LEDs_avalon_parallel_port_slave_chipselect      (mm_interconnect_0_green_leds_avalon_parallel_port_slave_chipselect),      //                                           .chipselect
		.HEX3_HEX0_avalon_parallel_port_slave_address          (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_address),          //       HEX3_HEX0_avalon_parallel_port_slave.address
		.HEX3_HEX0_avalon_parallel_port_slave_write            (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_write),            //                                           .write
		.HEX3_HEX0_avalon_parallel_port_slave_read             (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_read),             //                                           .read
		.HEX3_HEX0_avalon_parallel_port_slave_readdata         (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_readdata),         //                                           .readdata
		.HEX3_HEX0_avalon_parallel_port_slave_writedata        (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_writedata),        //                                           .writedata
		.HEX3_HEX0_avalon_parallel_port_slave_byteenable       (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_byteenable),       //                                           .byteenable
		.HEX3_HEX0_avalon_parallel_port_slave_chipselect       (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_chipselect),       //                                           .chipselect
		.Interval_timer_s1_address                             (mm_interconnect_0_interval_timer_s1_address),                             //                          Interval_timer_s1.address
		.Interval_timer_s1_write                               (mm_interconnect_0_interval_timer_s1_write),                               //                                           .write
		.Interval_timer_s1_readdata                            (mm_interconnect_0_interval_timer_s1_readdata),                            //                                           .readdata
		.Interval_timer_s1_writedata                           (mm_interconnect_0_interval_timer_s1_writedata),                           //                                           .writedata
		.Interval_timer_s1_chipselect                          (mm_interconnect_0_interval_timer_s1_chipselect),                          //                                           .chipselect
		.JTAG_UART_avalon_jtag_slave_address                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                   //                JTAG_UART_avalon_jtag_slave.address
		.JTAG_UART_avalon_jtag_slave_write                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                     //                                           .write
		.JTAG_UART_avalon_jtag_slave_read                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                      //                                           .read
		.JTAG_UART_avalon_jtag_slave_readdata                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),                  //                                           .readdata
		.JTAG_UART_avalon_jtag_slave_writedata                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),                 //                                           .writedata
		.JTAG_UART_avalon_jtag_slave_waitrequest               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),               //                                           .waitrequest
		.JTAG_UART_avalon_jtag_slave_chipselect                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),                //                                           .chipselect
		.Onchip_memory_s1_address                              (mm_interconnect_0_onchip_memory_s1_address),                              //                           Onchip_memory_s1.address
		.Onchip_memory_s1_write                                (mm_interconnect_0_onchip_memory_s1_write),                                //                                           .write
		.Onchip_memory_s1_readdata                             (mm_interconnect_0_onchip_memory_s1_readdata),                             //                                           .readdata
		.Onchip_memory_s1_writedata                            (mm_interconnect_0_onchip_memory_s1_writedata),                            //                                           .writedata
		.Onchip_memory_s1_byteenable                           (mm_interconnect_0_onchip_memory_s1_byteenable),                           //                                           .byteenable
		.Onchip_memory_s1_chipselect                           (mm_interconnect_0_onchip_memory_s1_chipselect),                           //                                           .chipselect
		.Onchip_memory_s1_clken                                (mm_interconnect_0_onchip_memory_s1_clken),                                //                                           .clken
		.Onchip_memory_s2_address                              (mm_interconnect_0_onchip_memory_s2_address),                              //                           Onchip_memory_s2.address
		.Onchip_memory_s2_write                                (mm_interconnect_0_onchip_memory_s2_write),                                //                                           .write
		.Onchip_memory_s2_readdata                             (mm_interconnect_0_onchip_memory_s2_readdata),                             //                                           .readdata
		.Onchip_memory_s2_writedata                            (mm_interconnect_0_onchip_memory_s2_writedata),                            //                                           .writedata
		.Onchip_memory_s2_byteenable                           (mm_interconnect_0_onchip_memory_s2_byteenable),                           //                                           .byteenable
		.Onchip_memory_s2_chipselect                           (mm_interconnect_0_onchip_memory_s2_chipselect),                           //                                           .chipselect
		.Onchip_memory_s2_clken                                (mm_interconnect_0_onchip_memory_s2_clken),                                //                                           .clken
		.Onchip_memory_SRAM_s1_address                         (mm_interconnect_0_onchip_memory_sram_s1_address),                         //                      Onchip_memory_SRAM_s1.address
		.Onchip_memory_SRAM_s1_write                           (mm_interconnect_0_onchip_memory_sram_s1_write),                           //                                           .write
		.Onchip_memory_SRAM_s1_readdata                        (mm_interconnect_0_onchip_memory_sram_s1_readdata),                        //                                           .readdata
		.Onchip_memory_SRAM_s1_writedata                       (mm_interconnect_0_onchip_memory_sram_s1_writedata),                       //                                           .writedata
		.Onchip_memory_SRAM_s1_byteenable                      (mm_interconnect_0_onchip_memory_sram_s1_byteenable),                      //                                           .byteenable
		.Onchip_memory_SRAM_s1_chipselect                      (mm_interconnect_0_onchip_memory_sram_s1_chipselect),                      //                                           .chipselect
		.Onchip_memory_SRAM_s1_clken                           (mm_interconnect_0_onchip_memory_sram_s1_clken),                           //                                           .clken
		.Onchip_memory_SRAM_s2_address                         (mm_interconnect_0_onchip_memory_sram_s2_address),                         //                      Onchip_memory_SRAM_s2.address
		.Onchip_memory_SRAM_s2_write                           (mm_interconnect_0_onchip_memory_sram_s2_write),                           //                                           .write
		.Onchip_memory_SRAM_s2_readdata                        (mm_interconnect_0_onchip_memory_sram_s2_readdata),                        //                                           .readdata
		.Onchip_memory_SRAM_s2_writedata                       (mm_interconnect_0_onchip_memory_sram_s2_writedata),                       //                                           .writedata
		.Onchip_memory_SRAM_s2_byteenable                      (mm_interconnect_0_onchip_memory_sram_s2_byteenable),                      //                                           .byteenable
		.Onchip_memory_SRAM_s2_chipselect                      (mm_interconnect_0_onchip_memory_sram_s2_chipselect),                      //                                           .chipselect
		.Onchip_memory_SRAM_s2_clken                           (mm_interconnect_0_onchip_memory_sram_s2_clken),                           //                                           .clken
		.Pushbuttons_avalon_parallel_port_slave_address        (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_address),        //     Pushbuttons_avalon_parallel_port_slave.address
		.Pushbuttons_avalon_parallel_port_slave_write          (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_write),          //                                           .write
		.Pushbuttons_avalon_parallel_port_slave_read           (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_read),           //                                           .read
		.Pushbuttons_avalon_parallel_port_slave_readdata       (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_readdata),       //                                           .readdata
		.Pushbuttons_avalon_parallel_port_slave_writedata      (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_writedata),      //                                           .writedata
		.Pushbuttons_avalon_parallel_port_slave_byteenable     (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_byteenable),     //                                           .byteenable
		.Pushbuttons_avalon_parallel_port_slave_chipselect     (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_chipselect),     //                                           .chipselect
		.sdram_s1_address                                      (mm_interconnect_0_sdram_s1_address),                                      //                                   sdram_s1.address
		.sdram_s1_write                                        (mm_interconnect_0_sdram_s1_write),                                        //                                           .write
		.sdram_s1_read                                         (mm_interconnect_0_sdram_s1_read),                                         //                                           .read
		.sdram_s1_readdata                                     (mm_interconnect_0_sdram_s1_readdata),                                     //                                           .readdata
		.sdram_s1_writedata                                    (mm_interconnect_0_sdram_s1_writedata),                                    //                                           .writedata
		.sdram_s1_byteenable                                   (mm_interconnect_0_sdram_s1_byteenable),                                   //                                           .byteenable
		.sdram_s1_readdatavalid                                (mm_interconnect_0_sdram_s1_readdatavalid),                                //                                           .readdatavalid
		.sdram_s1_waitrequest                                  (mm_interconnect_0_sdram_s1_waitrequest),                                  //                                           .waitrequest
		.sdram_s1_chipselect                                   (mm_interconnect_0_sdram_s1_chipselect),                                   //                                           .chipselect
		.Serial_port_avalon_rs232_slave_address                (mm_interconnect_0_serial_port_avalon_rs232_slave_address),                //             Serial_port_avalon_rs232_slave.address
		.Serial_port_avalon_rs232_slave_write                  (mm_interconnect_0_serial_port_avalon_rs232_slave_write),                  //                                           .write
		.Serial_port_avalon_rs232_slave_read                   (mm_interconnect_0_serial_port_avalon_rs232_slave_read),                   //                                           .read
		.Serial_port_avalon_rs232_slave_readdata               (mm_interconnect_0_serial_port_avalon_rs232_slave_readdata),               //                                           .readdata
		.Serial_port_avalon_rs232_slave_writedata              (mm_interconnect_0_serial_port_avalon_rs232_slave_writedata),              //                                           .writedata
		.Serial_port_avalon_rs232_slave_byteenable             (mm_interconnect_0_serial_port_avalon_rs232_slave_byteenable),             //                                           .byteenable
		.Serial_port_avalon_rs232_slave_chipselect             (mm_interconnect_0_serial_port_avalon_rs232_slave_chipselect),             //                                           .chipselect
		.Slider_switches_avalon_parallel_port_slave_address    (mm_interconnect_0_slider_switches_avalon_parallel_port_slave_address),    // Slider_switches_avalon_parallel_port_slave.address
		.Slider_switches_avalon_parallel_port_slave_write      (mm_interconnect_0_slider_switches_avalon_parallel_port_slave_write),      //                                           .write
		.Slider_switches_avalon_parallel_port_slave_read       (mm_interconnect_0_slider_switches_avalon_parallel_port_slave_read),       //                                           .read
		.Slider_switches_avalon_parallel_port_slave_readdata   (mm_interconnect_0_slider_switches_avalon_parallel_port_slave_readdata),   //                                           .readdata
		.Slider_switches_avalon_parallel_port_slave_writedata  (mm_interconnect_0_slider_switches_avalon_parallel_port_slave_writedata),  //                                           .writedata
		.Slider_switches_avalon_parallel_port_slave_byteenable (mm_interconnect_0_slider_switches_avalon_parallel_port_slave_byteenable), //                                           .byteenable
		.Slider_switches_avalon_parallel_port_slave_chipselect (mm_interconnect_0_slider_switches_avalon_parallel_port_slave_chipselect), //                                           .chipselect
		.sysid_control_slave_address                           (mm_interconnect_0_sysid_control_slave_address),                           //                        sysid_control_slave.address
		.sysid_control_slave_readdata                          (mm_interconnect_0_sysid_control_slave_readdata)                           //                                           .readdata
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clk),                            //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
